-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "7E4D7BEF6506AEEAFFB413DC32CFF16526FF02DA6DE6F26919551789DF1316D9";
    attribute INIT_01 of inst : label is "51E76ECC3B30298685794D6035B2249C04120535B24005C25FFDF24CB30738B0";
    attribute INIT_02 of inst : label is "870E38763578DB0C97498248C6493164AC018FBA55AD658F39249189790D685B";
    attribute INIT_03 of inst : label is "00000000000000000000000000001E3C0F8AA8841ACA8700A79904C8320F02A0";
    attribute INIT_04 of inst : label is "947FB28C954791EE6FFD800A0E30DC9469A470298D238B86AC1431D3AE1741B8";
    attribute INIT_05 of inst : label is "03291577F5064C60B5598282AD663A08397F777ADC8D36E59C9CA3C8F737FFCF";
    attribute INIT_06 of inst : label is "E626533270414A286A59000414D448393F5402C14028911188B1C6104B0FAC13";
    attribute INIT_07 of inst : label is "006B005E8E95D9DEC0DD6FAA3656B5083544E419871D458212880A9028DB16D8";
    attribute INIT_08 of inst : label is "B5963DAB6FA6C927FFAFF9E50B22264CB310005081A55414A062E1442EA0A47B";
    attribute INIT_09 of inst : label is "EC2FC5D80BA4D6A140B888C30466A8159328A2E08084D6B6230053719753B2B8";
    attribute INIT_0A of inst : label is "FFDFEC337F5B78D993FCF7FC67DE5D7F732832F13DB3E45A10D0BE67418560BF";
    attribute INIT_0B of inst : label is "3B999EB9939B34106829E8A00FDEA0829243F7BF9B692740FFC11F6686C800B8";
    attribute INIT_0C of inst : label is "00000001D3204744C32224001DC2224F770180E0380ECC3FB08D543032CC6B99";
    attribute INIT_0D of inst : label is "24CC6185C30266BCC679E6271E79E798F76DDC6F86170C0DDA29FB5A8B245223";
    attribute INIT_0E of inst : label is "61CF074667821381873C0C37030E06160C2700C2C06073781FF9FFCC3BBF5B6C";
    attribute INIT_0F of inst : label is "000000000000000000000000000000000000000099E284E1000041D199E284E1";
    attribute INIT_10 of inst : label is "09370744C3ED00011E32A798AF215801F6500AA108880F33808B0000D8C010EF";
    attribute INIT_11 of inst : label is "59AFCB10ACDA1800524E06E0E8AC3E9111119E59F91B2C8044120821BBFF8253";
    attribute INIT_12 of inst : label is "6331E98888A8AA080011964FAC8001454A00015BCDE4AAA0003BBE2530DFD600";
    attribute INIT_13 of inst : label is "0025DD902612402311589826C0733E4A334D9FE000143B88C54C66AF82B9891E";
    attribute INIT_14 of inst : label is "830279F70B2691007803069C96A0CC32942B68E053F97C74D3115CABFFFC8008";
    attribute INIT_15 of inst : label is "C9D00011151116532AB85A3311111189D409819137628111AC60882804D8100C";
    attribute INIT_16 of inst : label is "FE73FD2BA1D15E95D0968FFFC44443EA572150FA22A388D5620FFF0318982D2C";
    attribute INIT_17 of inst : label is "00C00544254256A822124496C925B49125B249247FFFF8705454547373E5EFD7";
    attribute INIT_18 of inst : label is "FB5DEC731911A2284588AB0727AC4094F9170D32CC500446C6001190B3A48248";
    attribute INIT_19 of inst : label is "0008099BF380E21A59C69844089CA2E189C48D18F000B26D48BB8C4AA02CBFD7";
    attribute INIT_1A of inst : label is "2F75761E01798009D96775761C02D361DC63111127D326DB2082659901293F9F";
    attribute INIT_1B of inst : label is "B3A2A161B613CF1EB062C24586488102DB640001095659976EC00F8008579AEF";
    attribute INIT_1C of inst : label is "00000000000000000000000000000000000000000000A00003F34E3300451899";
    attribute INIT_1D of inst : label is "D5A8080080008000203E8200240024002800400067A512007F80828A10068000";
    attribute INIT_1E of inst : label is "45A25547BD5479D5479CDE79F590CC96464BBF24BC9FA4D269349E0804AA9241";
    attribute INIT_1F of inst : label is "C7B06D1956DD5AA76E75E4263386642681805A00158186464924E2512492464B";
    attribute INIT_20 of inst : label is "00000000C62DC62DDC6CDC62A75F4744993E1080032695DD54F6E474D35D4A5F";
    attribute INIT_21 of inst : label is "80042803400007E69C7E008A31FF67465AC36C3340001B78E020361A00816D7E";
    attribute INIT_22 of inst : label is "96CB2CB297678A2028A6FC2E5000C100F055EE3250108BE2E09192000880D820";
    attribute INIT_23 of inst : label is "A2E08CF800AC9B14A5B8C4AA280B2FF5FED77B1CC645688B0B8181EBC4B23481";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000284C400C8099BF380E21A59C698440A9C";
    attribute INIT_25 of inst : label is "00000000000000000000000000000000000000018AA4470A9429349A42A0B618";
    attribute INIT_26 of inst : label is "E5170EEF800159362545862551A02DBFD7FB5DEC731B15A230B8607AF12C3480";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000032C04CDF9C0710D2CE34C22054";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "136116DD2700500500988018C11052400200118F7B46BEE1410A0B018E6313D8";
    attribute INIT_01 of inst : label is "1E54AC2080B278A252A37973903048B52E387290300801646D3EA2A00B22400D";
    attribute INIT_02 of inst : label is "C83441A11B0823203D7590E1A01EB38100A732A45C532CBB500E041DDEA701A6";
    attribute INIT_03 of inst : label is "0000000000000000000000000000587C9925C5A08A414E11EF881440B02F5062";
    attribute INIT_04 of inst : label is "A6AA853007792222D0080004380EED18B0E28161271403421DA74920DE0F0079";
    attribute INIT_05 of inst : label is "D42DA3FEF32290E4C1A61ED0F5A3392D098185FCD77E4A0A6001BC911168001C";
    attribute INIT_06 of inst : label is "C66BF116262D6EE5E4791495969DD98AC11CA6CE526CD22D91F8E2A15D457645";
    attribute INIT_07 of inst : label is "2C46B690C2315640C90EF6AE6D794B91C8880699943D699502CCD05C64373259";
    attribute INIT_08 of inst : label is "4AEA4740A1C00E037F5BFA22C68454200B22C97934128CF2F366E265BEE6948B";
    attribute INIT_09 of inst : label is "15484A20B0DD8AEA6969994E36086D2A2153942725498AEA7463AD9A244C8159";
    attribute INIT_0A of inst : label is "005411010125080101FDCBFD4920012E914A48B21556F83921C9151752330928";
    attribute INIT_0B of inst : label is "148A822A8163353310B451531496B1BD1490304002AA498000C9524B6A1B227D";
    attribute INIT_0C of inst : label is "000000018924CC21C30790000A00A0A0069381E048002F5803308A59802CA2AA";
    attribute INIT_0D of inst : label is "006CB2CA659489A6CB6DB648936DB6D902244C04DB29B6502AD64502E02B5670";
    attribute INIT_0E of inst : label is "078064B0B09C60CE1E06F0D1BC3B3B3E74C197478B862D8A3BFDFFD47C010102";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000002E2618330000192E2E261833";
    attribute INIT_10 of inst : label is "30D828589CB17333AB54D5A14B4293265AA99F14A5D11204D11D7ED7AD093460";
    attribute INIT_11 of inst : label is "EB4545BDF5A2AE4894007B050B29CB17333A84A6243F558888B538D00E9FA6A0";
    attribute INIT_12 of inst : label is "2C7ECF31111F34D1333AAAD6590888FB7BCE73A2D168AAA000042A4EC20A8B5A";
    attribute INIT_13 of inst : label is "914AA0214AA2A67473AD2140C92808D454922804CCA90199EEB10F4536D2D579";
    attribute INIT_14 of inst : label is "273DE483400C0595C8AE1EC169CC45105A6F6C4AA60A42BB6C23A1140152D394";
    attribute INIT_15 of inst : label is "6CF19187E3E3A5A4E65A920422223AC276521D23AEF0A53088E4BCA160592928";
    attribute INIT_16 of inst : label is "01843776EE9D7BBB775CB000088EACA6A53F3503CD15F3E8F45C800191673F3E";
    attribute INIT_17 of inst : label is "69C8B738B28B725907324496C925B49125B24925EAA80AA20899888B84063018";
    attribute INIT_18 of inst : label is "53254C9B2B3EA64217C2D338086916D2FA2596802C924A140E45840405E026AB";
    attribute INIT_19 of inst : label is "001F30ECB9ECC454CAF7A9231F09A45298C99A794971C1B5E4D5EE874CED85C9";
    attribute INIT_1A of inst : label is "082344B057963224804C2344B1270D6480F7B337F08137AEC715005A134A0040";
    attribute INIT_1B of inst : label is "0C44E66540138E9DE4C496892F245E64025B4D932520130522B644B225386040";
    attribute INIT_1C of inst : label is "00000000000000000000000000000000000000000000200002AAE85024C831A8";
    attribute INIT_1D of inst : label is "E6C008008000D555200B82003500240028004000745D1AD45D558293100A8000";
    attribute INIT_1E of inst : label is "ED7E088883998A0888A210964924103410188C0DF03981E0F07838F14D85B013";
    attribute INIT_1F of inst : label is "E30012926B1675EA8747D06B3556EA47307DA525299394101822E4D86034101A";
    attribute INIT_20 of inst : label is "0000004FD01CD01CECB6E0666E924048810A1280024343DC267C402C2F2B0261";
    attribute INIT_21 of inst : label is "6598791840000555D0A0499063501888CCCA808B520012F400203ECD018326C0";
    attribute INIT_22 of inst : label is "000240241D781064995AA8594964C931F24D6B046232B2A50612B024D19BDB32";
    attribute INIT_23 of inst : label is "A45215A4BB706C28735EE874533B617254C95326CACFA99914CC8A57CF51BD11";
    attribute INIT_24 of inst : label is "00000000000000000000000000000000DACC32DF30ECB9ECC454CAF7A9231F09";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000001A868A3019A2868341936F659";
    attribute INIT_26 of inst : label is "4D2296524B89E0DA730AF743A34CEC85C953254C9B293EA6594CB295F3D7BD11";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000016798765CF6622A657BD4918F8";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "00040400C20010010A340BD472DFE8AD007F00DC1691693068291C8E48A9D50C";
    attribute INIT_01 of inst : label is "9B76C844112438A210C3147600A08D213C38D700A01001F670BE82C61A422454";
    attribute INIT_02 of inst : label is "849C24EAF76B1245B05526C022DAA54DA529DB3614A5A8A3446C348AF74638FB";
    attribute INIT_03 of inst : label is "000000000000000000000000000042282BA1E1A003E04600EF880440300F5020";
    attribute INIT_04 of inst : label is "A6D585C80D2DB346DBF80008693568B957FC48208FE24097613A5A61A81400A1";
    attribute INIT_05 of inst : label is "D0202473B102D040F07F04707C230A03AD8257FF1F83FE2B940C96D9A36DF832";
    attribute INIT_06 of inst : label is "44313D9E2A294AB0D6519445149558EEB4C46A85502A900D00F8E3807145C4E1";
    attribute INIT_07 of inst : label is "034B90C400715C028851A62A82140282FCCC60D108590D084280B054A23A1D85";
    attribute INIT_08 of inst : label is "9FFE07FF6160AB01D56EABC0826EEDC61A048A1805A095703142215422A2843A";
    attribute INIT_09 of inst : label is "5C7BC89CE17D8EAB1A7939CD3528A148B37AA66F21CB8EAC7F63F6FAB1413243";
    attribute INIT_0A of inst : label is "7F0AA51420DB081501A96F556DFE0C3AD9CA16FB9F73AE1810C0863451A26A94";
    attribute INIT_0B of inst : label is "80EEC2FEE00AA7517C84FDF72EDE83BF96912255BBCB4BDE28856FEDEC5A32B5";
    attribute INIT_0C of inst : label is "0000000104E007A8E72D4000000AA004349481E05804414319ACD66A18682FEC";
    attribute INIT_0D of inst : label is "6C08020B0437C92080410408D041041030C184E0182C10DAD22FAE5AAB0E1E31";
    attribute INIT_0E of inst : label is "460002D4D43A601D1800E8D03A30342A6CC016A50B4616CF3AA7AA9E7F56386E";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000370E9807000000B7370E9807";
    attribute INIT_10 of inst : label is "B06CACC0D6D95273FA741F797EE2DA336EF19FC671FAA794911D9DC7FD585C4F";
    attribute INIT_11 of inst : label is "EBE3A25A75F2FA1526D96D95984D6DD5273FC6BB730D7D58C8FF2C91B5D523F0";
    attribute INIT_12 of inst : label is "C71BEBA1939DA69C363FBEFF7DC8D8ECA729CBF7BBDCE6C11B06967F594744B4";
    attribute INIT_13 of inst : label is "015BB0A14FB2EC7F73FD296298091CDF36DB9B60D8FD101B0FDCE3E1A0BAF90C";
    attribute INIT_14 of inst : label is "A20068A3416C3425712B940852C84518122240EAF4A14C6DB633F505DFBE10A5";
    attribute INIT_15 of inst : label is "8D6BB9A5B5F5F3B6C65E9B1433637FC2E678ADB1AAB0E141244081D1E010484D";
    attribute INIT_16 of inst : label is "C5D5D95B2BD91CBF97DE825F0D8FEFC2FEBD17A861879ACD66999FA989CF3636";
    attribute INIT_17 of inst : label is "088081588588001A81126596FB27B5F72DF77F2D95545EB29DCCCCDDD4E763DD";
    attribute INIT_18 of inst : label is "603180CA021F2842F15E1A492FE1FEE00F3FFA18694092D6548434B597E1AA48";
    attribute INIT_19 of inst : label is "00123037E046065803A5F8110F9FA2620C850B50F8DBE0DCE8F74BEFE2095F1C";
    attribute INIT_1A of inst : label is "F61243BC00D3A32837FA1242BD018740308532722230B7BBE5BE30D3B16F12BF";
    attribute INIT_1B of inst : label is "6EE78D41E300008150DE77FCEF421B29AA2D6591210DEA7B025463A3280D3618";
    attribute INIT_1C of inst : label is "00000000000000000000000000000000000000000000A00003C1D818204418CC";
    attribute INIT_1D of inst : label is "F8E008008000E666203C82003D44240028004000448813326E66828C10038000";
    attribute INIT_1E of inst : label is "0D262DDD8CDDD8DCCDAC42BB6DBC45B0D2DA8C6879B98DC6F371BC994501B0D1";
    attribute INIT_1F of inst : label is "C7071C921F4DB9BF2E336563EE824ECFD1010143490106D2D8A2E35361B0D2DA";
    attribute INIT_20 of inst : label is "00000049813D813DA9559272FA65464E891280848395652F847D16C5B7A9376D";
    attribute INIT_21 of inst : label is "6040398340000783B02040883110DDCC0A83C61A500000910040002000008200";
    attribute INIT_22 of inst : label is "924B6D921A800824086C546B40468110F144CF166130894629D0B020000890B0";
    attribute INIT_23 of inst : label is "A263117C6AF8362CF574BCFE188257C7180C603280874A18960C4BE687F12F89";
    attribute INIT_24 of inst : label is "00000000000000000000000000000000929682123037E046065803A5F8110E9F";
    attribute INIT_25 of inst : label is "00000000000000000000000000000000000000010585765623F371BCD124A490";
    attribute INIT_26 of inst : label is "F903121FC6D8F06EF58BA5E7F162085F1C603180CA001F28416082F9A1FD2F88";
    attribute INIT_27 of inst : label is "000000000000000000000000000000000000001E1181BF023032C01D2FC0807E";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "05AC0404420414410AA50DA893C920ED1028D885A27124B0501C02001C981208";
    attribute INIT_01 of inst : label is "BFBBCC4711F334020243949B0870660037BF77087008069FF023ADC517221480";
    attribute INIT_02 of inst : label is "82B415B0D1269F2DA083968236D0F24D2C66FDDE958180418068358A2B720DB5";
    attribute INIT_03 of inst : label is "00000000000000000000000000004A14ADA16301048046DCD080D826D9B0103B";
    attribute INIT_04 of inst : label is "1ED5918C0264B1C61A0B00082D0278581AE028221701400A8410010088046020";
    attribute INIT_05 of inst : label is "91C43089E32E4427E931A06769E2116BB6C0337D0D2B26635C093258E30D0403";
    attribute INIT_06 of inst : label is "5E61644213A4621C942AD2E0C70CE1742FC42A4B22A2674A9CC4014DA0068470";
    attribute INIT_07 of inst : label is "2292334606D12D29F1D42F4E52269018644450FCD5160AD0A8DE174E202127C0";
    attribute INIT_08 of inst : label is "D94E60C94363D300FF67FB10E3A27845173159018EC0E41202355220E4E618F3";
    attribute INIT_09 of inst : label is "5972A6EBD7BE8CD31A57FD2E3360A14A871E3BCC45988CEFE7BB3640D18DAA60";
    attribute INIT_0A of inst : label is "058BF610304A1C7A80FE2FFC2CB18A10FCD45A4B8A610D5A5AD29E27A2ABA9D7";
    attribute INIT_0B of inst : label is "91A88DF461839A33C999CB27A24E1F39A621A74498C3021FA84C292E8E52AA50";
    attribute INIT_0C of inst : label is "00000007C3C40C868E0000001FEAA0462EE380A00802ED01B596C961145CDF44";
    attribute INIT_0D of inst : label is "2754EB8B5536E455CEFBAB662AFAEEA99A5CAA5FAA2F545CD06DBAD0FAEE6871";
    attribute INIT_0E of inst : label is "7641027E7FBB719DD905EEF17BBAFDBAFAE333B739F6066D5153FFCAAA929725";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000009DEEDC670000409D9DEEDC67";
    attribute INIT_10 of inst : label is "3864EC0A4E7C2FBF3A6213BF6772C8873C39FBBDAF9ABB30F5FAD696B0714059";
    attribute INIT_11 of inst : label is "D960A7096CB0385586486C8D8104E7C2FBF3E33193BB18BEBFD68E14905FC73C";
    attribute INIT_12 of inst : label is "D2F72CB37DFBA69EEBF38C5965DBAFDDAD394F39DCEC50514167157014414E52";
    attribute INIT_13 of inst : label is "1983BD8D8E34CFE7AB300D62F11B46C72659D13BAFCE18757CCECE60C6CA9C34";
    attribute INIT_14 of inst : label is "A12948210368348C3C618E5A408020101221A52234B14545962F3C256A0E10A4";
    attribute INIT_15 of inst : label is "B145FD81717137B3952C0D31FFEAF30087DAA6B98AB14479642628D1A009082D";
    attribute INIT_16 of inst : label is "74F06B3D673A359EB3B91A55BAFCF646327631A86186994CA64515CFCD89E460";
    attribute INIT_17 of inst : label is "08CDB91C91D98219003244B6E965FFFFBFB77FBE155754334444445470B9F2A5";
    attribute INIT_18 of inst : label is "24B490D92A998DE8F99F1131253ABBE1073A78145C8042DA426DB5B5B2A1A361";
    attribute INIT_19 of inst : label is "0014B83275546FC90B20B913CCE58522CA494B6928CBB0CCC7F740D6625512ED";
    attribute INIT_1A of inst : label is "266B86E033570AA699262B86A1668F269AD7BEAB539BBAB5D7D628BBD3771AF5";
    attribute INIT_1B of inst : label is "AAA7DEE4E2A4512249A2DCC5BA226FACCC6914132426499270D11C8AA535734D";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000020000280CA0D24441166";
    attribute INIT_1D of inst : label is "8118080082AAF87820008A003EAB24002800400045181E0E7878829F100C8000";
    attribute INIT_1E of inst : label is "58040555254450444504C60B2CB055A0D6D0266AD1A8CD46B351AC11280110D1";
    attribute INIT_1F of inst : label is "45613453034438BAAE990220A41A4846194B49010C9096D6D041159B41A4D6D2";
    attribute INIT_20 of inst : label is "00000061851A851AB81A8A42630D4140812A0004928101045CDE301625B5723D";
    attribute INIT_21 of inst : label is "644F339A40000501940A48882245554CADC9C513A20000100000090000009000";
    attribute INIT_22 of inst : label is "96D92492100088A5A865576B9C55CA2C0388E497F8B715762DC3194418486979";
    attribute INIT_23 of inst : label is "0727551462EC32AE63740D67189544BB492D24364AA6E37516BA8B23CA710589";
    attribute INIT_24 of inst : label is "00000000000000000000000000000002034C8014B83275546FC90B20B912CDA5";
    attribute INIT_25 of inst : label is "000000000000000000000000000000000000000102020A08043349A0D580B279";
    attribute INIT_26 of inst : label is "2C2916194669D86463ABA06B39625412ED24B490D928998DD16BA2C8F29D0589";
    attribute INIT_27 of inst : label is "000000000000000000000000000000000000002225C193AAA37E485905C89E65";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "04202090C20353354B4945058082480A142A556086C9050460204822000D8C01";
    attribute INIT_01 of inst : label is "8B66E845112778806280B7574A2ACE8A725EFF4A2A180197F2038AC51267528A";
    attribute INIT_02 of inst : label is "CA4652311A0026602689309ED011266101CDDBB68801A0C281098430633A1BBB";
    attribute INIT_03 of inst : label is "000000000000000000000000000040C990350DC9440D4655F70C5442A8AF394A";
    attribute INIT_04 of inst : label is "E6D5808841E5B3441B5F80042C894121A09CA549C4E52B6312084200D2090148";
    attribute INIT_05 of inst : label is "B9A4A202933D598DFCB92FED68E601474DA9560419012E215448F2D9A20DAA92";
    attribute INIT_06 of inst : label is "144FA6781A252458A43D90A49288E3414809A49A6646522815E08345610182F3";
    attribute INIT_07 of inst : label is "6665320403F71C209306B9245B2048514CED568016A26813BA46564F54A82066";
    attribute INIT_08 of inst : label is "A3CC4DDBA777CB21D46EA3B2E46676C5126239231D1288A647061274AA6C9588";
    attribute INIT_09 of inst : label is "5962B911DA030E4B3B7B9BDC70E4C7696418B094ACFC0E4DE6FF3242814A5B41";
    attribute INIT_0A of inst : label is "456BE85224DD3EF990A86D526DB58EB2C66CD6DB5B7B2F696B5900246688A354";
    attribute INIT_0B of inst : label is "001111013882A662DC939A6EB6D89319D6450E4DB2EB2A1F291AAB6C0442EE61";
    attribute INIT_0C of inst : label is "00000007082C05288A7AAA000AA00E8424A681A04800BB6125B2DB6314499013";
    attribute INIT_0D of inst : label is "6CA88A2B96564038081104421C41441134C182C82CAE51D982C01082504098E5";
    attribute INIT_0E of inst : label is "0E4A6CE8E850F2283929C1F67070A86951E6590D6C8E424FA402AA8F0A36B06D";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000003A143C8A00001B3A3A143C8A";
    attribute INIT_10 of inst : label is "7927EF5AEEF973373C72D7356E6ADEC77E3FFBE73B9996F3FF7A318E31533034";
    attribute INIT_11 of inst : label is "D871F0BCEC32304CC6DEE4FDEB8FEF973373B6BE3E2A1C8889D7B6D5BCF5453F";
    attribute INIT_12 of inst : label is "9C536DB71179B6DA22730E5B6DBCCFCF7BCE773399CCAAF2ABC6D470D663E139";
    attribute INIT_13 of inst : label is "B72333972CBAFFE6EF30AF6A139F2D8656C9AD2889CC5C119CF78A7184D99D6F";
    attribute INIT_14 of inst : label is "2C648002900885B4B5A50CC140D044034ACE4D7038BE56AD93FF3C956B9E56B5";
    attribute INIT_15 of inst : label is "1E6919833373341351109B7337227302CBDA972BA890CD28C98C9DD3A603AB60";
    attribute INIT_16 of inst : label is "57335F1BE3993F9FF3DE9395089CF8E637BD31A9659799CCE649950DE9C9F677";
    attribute INIT_17 of inst : label is "2B1A926D97C925532C7244B6C965B4D92DB37DBF955558870CCCCCDD32BCFAB1";
    attribute INIT_18 of inst : label is "663998C236BE275632C6527909531A730BB6581449E6EA1C18D4840401083529";
    attribute INIT_19 of inst : label is "00367912E0DC9D5D03A43932DF6FA57ED19F53D379F7B248877648CE667B370E";
    attribute INIT_1A of inst : label is "6E03550A93938EA4336643554BA7064C30C72333B7321CB35DD62897166B12C5";
    attribute INIT_1B of inst : label is "66675A5562EC30E14B8680CD02266BA59A529256AD2CDD3606A9820AA739361A";
    attribute INIT_1C of inst : label is "00000000000000000000000000000000000000000000E00002A308EF24846B57";
    attribute INIT_1D of inst : label is "D5CC0D57F199FF802A6286113F6D36693D5573334C1A1FFF48FFAAAA1116F998";
    attribute INIT_1E of inst : label is "B8DC7CCD36CCD36CCD15CE5B6DB154221013370F542EA150B85C2E510C158816";
    attribute INIT_1F of inst : label is "35F202506C1AC2C28165A10A396384001825256DAC363010114C85484C261031";
    attribute INIT_20 of inst : label is "00000065B482B482C1A0E93403BB7F7EFDF3B70CB210424483510C2995024501";
    attribute INIT_21 of inst : label is "60CB7789C000054611C64908D662CCCCACAAC512660004000010000000400000";
    attribute INIT_22 of inst : label is "BA69A6921500084C9027546B4D548D3D024ECC17EA229D66A452804C205991BA";
    attribute INIT_23 of inst : label is "257F573CFFEC92EC63648EE7599ECDC3998E66308DAF09DE562A2B728E712198";
    attribute INIT_24 of inst : label is "000000000000000000000000000000016A1802367912E0DC9D5D03A43933DE2F";
    attribute INIT_25 of inst : label is "00000000000000000000000000000000000000016C49CAD138B044261D5A40C1";
    attribute INIT_26 of inst : label is "793BF51BCFAFD92463AB24773A667A370E663998C234BC2765628ADCA39D2199";
    attribute INIT_27 of inst : label is "000000000000000000000000000000000000001133C89706E4EAE81D21C99EF1";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "6800200042035335374091248000590B00F455E48248248000400002000B0009";
    attribute INIT_01 of inst : label is "AA5EB8C83243751672895C532140481EF89D6F21400D5135FE42168824230000";
    attribute INIT_02 of inst : label is "C006002010000A20345210C4A01A430380A552F41C124145890C0418521B52AA";
    attribute INIT_03 of inst : label is "000000000000000000000000000000409975454498454F55D09552AA92A0136A";
    attribute INIT_04 of inst : label is "CEAAC0291521A34C149F800008004000008001080400080200000200C0000100";
    attribute INIT_05 of inst : label is "1324A2894223C087E4AA1D7F5881C1254DA416855B424320551890D1A60A4A54";
    attribute INIT_06 of inst : label is "2868F14243A5667AA53FD68CB288914A088CA60A5266522A55C51515228C8F60";
    attribute INIT_07 of inst : label is "26F7728C4A789C8509063B645B2848D1CECCE2E650B92A5026C0594D74A2A15C";
    attribute INIT_08 of inst : label is "026855DB60629B45D56EAB42866664CC342269211D52AC9242D78AEC80459484";
    attribute INIT_09 of inst : label is "93450803F004AE63397FFF0EB200672C105294340468AE4974ABA48123485141";
    attribute INIT_0A of inst : label is "DE5E203048DB0453A2A84D544D3219BAD54A76FB5F6BAE73639B4478D38061A8";
    attribute INIT_0B of inst : label is "E2AAA10A869C45235F90986E16DD9FDDF603324DB6DB06205D0D3368009AAE58";
    attribute INIT_0C of inst : label is "0000000508A4CC00088000000AAEBE88481380200800A55E25329943209090A8";
    attribute INIT_0D of inst : label is "6D98CF2B9E5640792CC249423CD3092534D9B0D13CEC7959A6D0140640801463";
    attribute INIT_0E of inst : label is "979622606114652A5E59D2DA74BCE2BDC2C05057A816B6C116A6AABA2636366C";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000001845194A000008981845194A";
    attribute INIT_10 of inst : label is "306D2D4CCEFB2EEBB27657376E6ED80F7EB75F8C61D99210B75F18C730C921C0";
    attribute INIT_11 of inst : label is "F261E05AF93EBA4C86DA6DA5A90CEFF2EEBB5638386E59FFFEE61859B4F525B1";
    attribute INIT_12 of inst : label is "00DB659FFFDD9658EEBB2C9B6DBBBAEC6318C3B399CCFFA3FE84A9586083C0B5";
    attribute INIT_13 of inst : label is "9D03200508369D74BBA0116609080F96B01B5BD3BAE820770EC01B618C5BDB2E";
    attribute INIT_14 of inst : label is "2424F1C5880C0494F0A74C414934A8B35A664672B1C5696036EBA016D69E7294";
    attribute INIT_15 of inst : label is "68F777B7A7E7A024E64C5B90EAFFBB09A65B940BACD6A52208859EE7E0E1A920";
    attribute INIT_16 of inst : label is "88009652CA7B7B3B6739B4BA3BAE80ACA5F5655B6DB69349A4C36EF1D9B93FBC";
    attribute INIT_17 of inst : label is "290B9B2F93F9A95127336596FFB7FFB7F7FECB64BFA8B46B0CCCCCF491D2774B";
    attribute INIT_18 of inst : label is "60B182E622BA65C23BC7543E4AAC7E66FA74D12090826A10885C850504A43639";
    attribute INIT_19 of inst : label is "0016B2B6E6451D58332D31765D0D666EDB0D5B4169F564DEA7665AF76EE9372C";
    attribute INIT_1A of inst : label is "4C8B6033F6AA8AE432648B40732D548533856AAA3736592255144123D26B370B";
    attribute INIT_1B of inst : label is "44444295445BAE5CA39626AC4F264A259A00C153256CD936820C508EE56BA61A";
    attribute INIT_1C of inst : label is "00000000000000000000000000000000000000000000A00000800075A4C939AA";
    attribute INIT_1D of inst : label is "E6340B35FF8780003FDBFE3C3FD63D332CE64F3C544817555DAA9A93104A981E";
    attribute INIT_1E of inst : label is "7E3F0ECFECCCFECECFEE021A69A0E838101ECA09E8350180C060345568355A13";
    attribute INIT_1F of inst : label is "01F0001000000082000100002002000012252525AE1210101C3196487838101C";
    attribute INIT_20 of inst : label is "00000045B000B0008000800002007C78F1E3B629020000040010000001000001";
    attribute INIT_21 of inst : label is "64CD75914000010000F3499273D8888B952A8824520000000000000000000000";
    attribute INIT_22 of inst : label is "09009001140016E5B94AA954DD4D0B6502DD48A56AF2BA9546761AA4D1D9017A";
    attribute INIT_23 of inst : label is "E66F5534FA5937EF5265AD775BBA4DCB182C60B988AE197057393B768B6169BA";
    attribute INIT_24 of inst : label is "000000000000000000000000000000016A8C0816B2B6E6451D58332D31765C4D";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000001600002C00010703C195A6C55";
    attribute INIT_26 of inst : label is "6F33761B4FAAB26F52AB2D6BBB6EE8372C60B182E620BA65C573CEDDA2D969BB";
    attribute INIT_27 of inst : label is "00000000000000000000000000000000000000023595B73228EAC199698BB2EA";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "364912CB61070F70FF66619E16DB646D127F4476D96DB6F9717E19099FD99D94";
    attribute INIT_01 of inst : label is "0B60EE6499392C91386114BF843D240A3C1CE7843C2665A73322A0E49382FFF8";
    attribute INIT_02 of inst : label is "BFC5FE3F1FF8918DD451C75486EA394E2E319B06E1C824D2A46539C36B6E08BB";
    attribute INIT_03 of inst : label is "0000000000000000000000000000173E45D0709A40C43644B74C4662288F0908";
    attribute INIT_04 of inst : label is "A6D5C1B0660DB1661FF87FFF8FFC7FFFF8FFFEF7C7FFF7E3F8410410BFFFFEF8";
    attribute INIT_05 of inst : label is "095218039993C6327639C0E05E213C907AFD96859B7B6F23246B06D8B30FFFDA";
    attribute INIT_06 of inst : label is "872211119B329108948CBE0201265C3A2EE211E399112981CCA493446933A2E1";
    attribute INIT_07 of inst : label is "98313C77865B6610EC9CED13B6CF22CE0647695DC58991C421390065120785C0";
    attribute INIT_08 of inst : label is "91AF39DBC1720301AA6D53CC19232064939C9ECEE9CC632D9C72C8231F326B1B";
    attribute INIT_09 of inst : label is "D863C4C9F9650D2B942311EC3C231284D75B424539890D2E5732B6E69DB16408";
    attribute INIT_0A of inst : label is "7FCAA4D1BEDE0E4081556EA96DBE4D30F11332C318630C8C8464373719806497";
    attribute INIT_0B of inst : label is "B9888C9AA3C339990DCC882646D8411D860DD32DB0C31A40FFE56B6D8D486323";
    attribute INIT_0C of inst : label is "00000004E2D227FE10D002000AB441672658FE3F8FE2E187B0C06024924E49AA";
    attribute INIT_0D of inst : label is "24CE278B4F16E41CE679E7260E79E79C9E4C984E9A2D345DB11B72110263E72D";
    attribute INIT_0E of inst : label is "4605966666D7608B1814D8D936326C28D8C915850AC616FB2957557E57B21324";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000009BB4D8220000659B9BB4D822";
    attribute INIT_10 of inst : label is "B26CACA0DEFC8222BB6707B36D62DA277CB11794A55C4B9051165295B36C920B";
    attribute INIT_11 of inst : label is "BF6D8F6B5DB0BB2216496D9D942DEF88222BD6B9B13F5DCCCCB6410892CAB3B0";
    attribute INIT_12 of inst : label is "426B71C11115C718222BAEDB6D8888ADAD6B5ABB5DECAAA000379439115B1ED6";
    attribute INIT_13 of inst : label is "494BBC814EB0C45622B06D7BEC710C5666DB37E088ACDB116ACC4D6DA71A588C";
    attribute INIT_14 of inst : label is "93921C7233643A420210271C241064892111F26AB3FBDCCDB622B443FE592842";
    attribute INIT_15 of inst : label is "894111C8B8F8B6372231AD9022222B069B5EC1B94AB932932E704DC1E31C848D";
    attribute INIT_16 of inst : label is "FE51DB5B6B9C9DBFB79E4E7F888AC2D2B63695FC71C64C2613015F034C892424";
    attribute INIT_17 of inst : label is "84E0C8C5CC5C870C93924496C925B49125B249245557F9834444447651E17787";
    attribute INIT_18 of inst : label is "603D80F3999310E8E89D03976FE4D7FA0BF69E924E1920E6E70639B9B719D064";
    attribute INIT_19 of inst : label is "000C3036F300EE581B81BC8949CC9266C1E4C33C648160D8B03702E5712CB68F";
    attribute INIT_1A of inst : label is "2C63B61E0843A633996C63B65ED086739D9DA322D6931DBB05D7249B99739F9F";
    attribute INIT_1B of inst : label is "22328472724861C340E2C2C587912BB0DD64801DFA865B967CC80FA6328433CF";
    attribute INIT_1C of inst : label is "00000000000000000000000000000000000000000000FFFFF8FFE33132308C88";
    attribute INIT_1D of inst : label is "F9FC08F6F87F800020FC9E6024C63EFF3C0740C0458516336ECC878C11D3F9E0";
    attribute INIT_1E of inst : label is "D4620467AC667AC667AE421B6DB355D4E6E88A6429914CA643A1D503E69088E8";
    attribute INIT_1F of inst : label is "F10FFF1FFFFFF8E3FFF1FFFE3FE3FFFF1390909085C9C6E6CA281083A1D0E6C8";
    attribute INIT_20 of inst : label is "00000050CFF8CFF8FFF8FFFFE3FC40408102480927FFFFC7FF1FFFFFF1FFFFFF";
    attribute INIT_21 of inst : label is "7B3121E3FFFFF1FFC66A64611914446508E4E493980000000000000000000000";
    attribute INIT_22 of inst : label is "600092481000E11E466E542A2480E0840824AC97582D4942B18988332E4E7E39";
    attribute INIT_23 of inst : label is "926614B24158362C59702E571C4B2DA3D80F603CE664443116998B6565700DC4";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000321E5060C3036F300EE581B81BC8948CC";
    attribute INIT_25 of inst : label is "00000000000000000000000000000000000000019FFFE33FFE0B29D0E8C9073C";
    attribute INIT_26 of inst : label is "649334DB2408B06C590B8172B8712DB68F603D80F39B9110D169E2D959DC0DC4";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000030E181B7980772C0DC0DE44A46";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "3249364B61060E60FF2C008C32CB206F407F00C2CB24B2410101010340584098";
    attribute INIT_01 of inst : label is "0924444411102882304104CA0010240038184600100784A32000024411020000";
    attribute INIT_02 of inst : label is "8004002010009B04D4508354826A114624208922C48030C38035188B39780899";
    attribute INIT_03 of inst : label is "0000000000000000000000000000163C0DC0208001C01600B7880440300F0020";
    attribute INIT_04 of inst : label is "2655C0B0078491444FF800000800400000800000040000020000000080000000";
    attribute INIT_05 of inst : label is "0160518D40118462D41B804450011000337C92808A2927212409C248A227FFDA";
    attribute INIT_06 of inst : label is "022115120A23020094113C0411C010382EC40341D020310088A0820041870641";
    attribute INIT_07 of inst : label is "006330C60659300068908020000E02880644614C811D0080022C0A4420050DC0";
    attribute INIT_08 of inst : label is "91243C8960220900AA2551E04323644411109808888044201022404434008C19";
    attribute INIT_09 of inst : label is "C92BC4C9EB210609100311A82122220492CB86C5A08D060453229260B1C32018";
    attribute INIT_0A of inst : label is "7FCAAC103E4B0041005524A9249F0D16755A3251092164120082162251806097";
    attribute INIT_0B of inst : label is "91888D9881011D010D8C8826024C811C9201F32492490240FFC4492484446230";
    attribute INIT_0C of inst : label is "00000005C2E00400000000000AA10046225180200802E007B180C06010445988";
    attribute INIT_0D of inst : label is "24446799CF12642C4638E2241638E3889A4488479E673C4C9209263206237421";
    attribute INIT_0E of inst : label is "44074AC6C7D7418B101CD89B36266C20D88315840AC412733554557265921124";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000B1F4D062000052B1B1F4D062";
    attribute INIT_10 of inst : label is "A024A4C05A690222913C039327264A2537911694A5480990D114569510681159";
    attribute INIT_11 of inst : label is "A624C529531392001249449C9825A690222952999914CB4CCCA20808926AA190";
    attribute INIT_12 of inst : label is "422920811114820822296589248888A4A5294A99CCE400000033947910498A52";
    attribute INIT_13 of inst : label is "09691C816492445222900D236839063232491FE088A419112A4C4524A20F4906";
    attribute INIT_14 of inst : label is "C30048230134180800000208000044100023A22F97F91C6492229403FEC82000";
    attribute INIT_15 of inst : label is "8141110090D0921322383690222229009B4880917105A3136C608481C0080004";
    attribute INIT_16 of inst : label is "FED1CCC999191676CE988E7F888A466193370CF82082582C16051F034D882420";
    attribute INIT_17 of inst : label is "10C081058058020003124496C925B49125B249245557F8224444447651F177C7";
    attribute INIT_18 of inst : label is "3214C851191320E8618C01176FA5D54A01A2881044100062460419999720C2E8";
    attribute INIT_19 of inst : label is "000C201271006E4C8905104509C4A2270144812820814048A0620A4528AC9385";
    attribute INIT_1A of inst : label is "2422F20E14C1E622992822F24EE98222999CE2226391111104D2208910391F9F";
    attribute INIT_1B of inst : label is "223600232248614201224044810029A0CF248030E3464A923E480766234C134F";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000020000080023160501888";
    attribute INIT_1D of inst : label is "81CF0808FFFFFFFF20C083AA24383FFF2BF8400065011A0F78F0FEFF1E3C8600";
    attribute INIT_1E of inst : label is "552286478C6478C6478E4209249044D062688A3228D546A351A8D003C4009061";
    attribute INIT_1F of inst : label is "0100001000000082000100002002000013000000048182626A2880C1A8D4624A";
    attribute INIT_20 of inst : label is "00000040800080008000800002004040810200124A0000040010000001000001";
    attribute INIT_21 of inst : label is "4910212240000100046AC0A03154446D08464411D00000000000000000000000";
    attribute INIT_22 of inst : label is "492400001000A4B52A26546A500041400054A4135025A946A09590212A02EA31";
    attribute INIT_23 of inst : label is "A2263890415012245020A4520A2B24E14C8532144644483333998935412028A2";
    attribute INIT_24 of inst : label is "000000000000000000000000000000020140000C201271006E4C8905104508C4";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000001000002000009A0D068802228";
    attribute INIT_26 of inst : label is "251138490408A024501905229028AC93853214C851191120F339E24D50C828A2";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000032610093880372644828822846";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
