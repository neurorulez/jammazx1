-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "20E20E278EB80406894E2E0E3E3838FC577D55555555555555558C30EB4DF389";
    attribute INIT_01 of inst : label is "978E0896278038025F2690304ECD2FCED4538E4E13FDD7838BD75E20BC2A224F";
    attribute INIT_02 of inst : label is "AE0E1777771419777F57174014D8D09050A381E3B81E3A38078D7FCE384E01E3";
    attribute INIT_03 of inst : label is "E2A2F018BE26AEAE99F8E23E0E2DF88CE3E23884BE5C2F89F838B7E00E35BE7C";
    attribute INIT_04 of inst : label is "A9AA5550A63AA86F0AFE9BAB683AAB86AB1E63B1BA23FAAF188D28BD222F088B";
    attribute INIT_05 of inst : label is "D440BABAAD440EBE5502F7EED540EBAB6AFB55200BA6AEE02E9550FEEAFA039E";
    attribute INIT_06 of inst : label is "FE0AA9EAFAE0BAF7B7AF560150302BBEBAB80BE6A1FB72F80BE5103AAB5103AA";
    attribute INIT_07 of inst : label is "AFA021E6AC08557B01C0601C0601807022F7EEE002A0682AB6A9BFAC2FD55555";
    attribute INIT_08 of inst : label is "DBD50EAADAFBE9580FBDAAB80069AAE00AADFB802AB5543EF6AB805A01608FBD";
    attribute INIT_09 of inst : label is "88B679D26399E6F99E679AE5CFE30DB8AD2A2528F4FFE3CAD280482EEC0ABBBB";
    attribute INIT_0A of inst : label is "AE2E7F1FC2F03D84B6288AAF31E3C2F4A8BC2E2F8B8BE222F08870EF747F3C2F";
    attribute INIT_0B of inst : label is "6F4514B61544776AA7E7709072E685AECBE78B9A26BB2D6ED23EBEE2FB8BFEE1";
    attribute INIT_0C of inst : label is "E9F9F9CB02E033F8BCF7882D6682EE2DD262A7E7BDE2A1AFE2A1A38A863688AE";
    attribute INIT_0D of inst : label is "9A04B8607F23E3C3F8F0364BE1B4BD222FCB8BC062F898BC222F88ABA9D8E2F3";
    attribute INIT_0E of inst : label is "A22C611E334FCD7CE0BABC3ECE989BCBABC8BD222F09ABBB9F9CAF4A06224B8E";
    attribute INIT_0F of inst : label is "888888888A8AAAAAAAAAA888A8AAAFFCE7E707DA592EA6222F8A1EB5BC8887BC";
    attribute INIT_10 of inst : label is "AAAAAAAAAA888A888888888A8AAAAAAAAAA888A888888888A8AAAAAAAAAA888A";
    attribute INIT_11 of inst : label is "8DAB88888888A8AAAAAAAAAA888A888888888A8AAAAAAAAAA888A888888888A8";
    attribute INIT_12 of inst : label is "8833D2D20B4925931B4810F2AAD34F18FD2DDF8EABCBE31C32F8EF67AE1E9688";
    attribute INIT_13 of inst : label is "97C5FFD5A1974A51E116AD1B46A08221F254FB4EE33F4F4F0F15FDD6206B7775";
    attribute INIT_14 of inst : label is "C8BF88F89F0BF0AF0BF0AF08F0AFC9FB55965561ED954F0ED6AA61A553C3B6AA";
    attribute INIT_15 of inst : label is "AAFADE7763E7AAFE5920798BD9EB03CC07B60F19E7FBFB222678E0F3F458822B";
    attribute INIT_16 of inst : label is "F9EAABC60F3F72183C67E7AAEA28F35B3B91D7DA1183C54ECA062D23EA0AF3A7";
    attribute INIT_17 of inst : label is "512825B59DEEFE7AAEA0F39CD8E7AF19EF83CC87360F1F9EAABDFE7AAE90F3B3";
    attribute INIT_18 of inst : label is "626E74E742A2A2A2A2AE889E027809E3278CBC12FD67FDC0029000814FDC7B9E";
    attribute INIT_19 of inst : label is "3A1E8F2893C4C3B434D0040C6100B7C8FAD218CF2880988E74E74E74C888E74A";
    attribute INIT_1A of inst : label is "CBC062F82A0A92F02F00838C72F838BC02E00C3C38986B098219A999B831E8F0";
    attribute INIT_1B of inst : label is "942425E2CD2E79BE7499D38E17D3D39F55F695F470C3A39C2D9F126A22AB0B88";
    attribute INIT_1C of inst : label is "8B81E074EDA3B708C357FAFD4F5D4BB4077D5E38D4F5CAA3AAFD4F5D4B406198";
    attribute INIT_1D of inst : label is "C2023489F3002F00F8C0683818B7A2C4F0B2BC1F88C2327CCFDB4AE07382EAC3";
    attribute INIT_1E of inst : label is "227C2C0D2A7C2C882CE068184B38780A24E4B38603B00F00F02CAD22702CE818";
    attribute INIT_1F of inst : label is "4BD28BD07803C2192FA84BEA12FA84BEA2F2B88F38F38431F8878E1AF8C1E20C";
    attribute INIT_20 of inst : label is "A8A8A8AAEA68E8A8E8286868A82828286A2AEAEA6AAAEA8FC0B8C00F0AAAABE2";
    attribute INIT_21 of inst : label is "5555055D55055D550D924655D51951D185575504545054546595955154455568";
    attribute INIT_22 of inst : label is "24455D51951755615715415755615755615755635491506544541D55055C5585";
    attribute INIT_23 of inst : label is "7D8FEEBFD1955855455455C55C55855C50C544559559558514558555555554D1";
    attribute INIT_24 of inst : label is "15415655655635491506444543E09DFB62EDA9EF8D168AF96F97B7B868F8403D";
    attribute INIT_25 of inst : label is "9D924655D519151DC45155555554155155157156157156145156155555555145";
    attribute INIT_26 of inst : label is "5555555555555555D55555555D55551151D51951151D51951151D51951151D51";
    attribute INIT_27 of inst : label is "1864B05DD34F1C3310C3DD2495D5416554545511014555554554555554555555";
    attribute INIT_28 of inst : label is "BAE39EF8EB6EAB92A57E3CD0F05FDABC785AB7783861AB8F3C8F206AFB01ABEC";
    attribute INIT_29 of inst : label is "DBF9D45F945B0EA51EF3BD26F6FD1B8EA47BCEF49BDBF81B0EA9D1EF49BDFD8E";
    attribute INIT_2A of inst : label is "7C9663EC3AE5CEE3AAA56FD20AC3A947BCEF49BDBEBAD17BCEF606C3A91EF49B";
    attribute INIT_2B of inst : label is "E69BB7A8B779EB8B8E946AE709E9AC7CEA73B8EABC5BF454F0F081A77A3EC3AE";
    attribute INIT_2C of inst : label is "1B8EA9D30683AAFC798388385F6AAAAAAAAAAA8B7512D7F2EEEEE97F2CBBA2ED";
    attribute INIT_2D of inst : label is "A6EB8A9BAF145B4F26EEBAA1D3F78B3BDBDD1C46E3AAF7DE22343384DAA20488";
    attribute INIT_2E of inst : label is "AD0AAADB34ADA26BEF2E2D3889BB7673C9D1820D03AFD2689FB0A777B749BAC2";
    attribute INIT_2F of inst : label is "F8887AC322F088BC262F8B8FE0F02EAD0BE2AD073CAF80C3B8DA1ABEA2D2B698";
    attribute INIT_30 of inst : label is "F89DB9AF4BE3F8D0E7466D6F34BE222740FE39AF4BF829ECD236D22BD00BF222";
    attribute INIT_31 of inst : label is "F874089D30D334AF42F42AE210E23D223E3FCAF8D34089D27B234A3F8AB234A3";
    attribute INIT_32 of inst : label is "2274E1DF48E0AF42F42AE210F2BE37874BE262F0183E30778639EC8D2AB234A3";
    attribute INIT_33 of inst : label is "8D89BEEA1A26A274AE589BC6BAFCBE76AD2AD2F4E3488934E274DD3F4E23889F";
    attribute INIT_34 of inst : label is "AC26AEB89ABAF2ADDD2061884AE9884AE9884AE9884AEFB46E1DE3A8BEEABAAA";
    attribute INIT_35 of inst : label is "E22787AE23889E3C0B78E23F6CB73BB705A8BDC376A2F88F34BC061C30E7EDD3";
    attribute INIT_36 of inst : label is "F505EF7BB503BEEC2FFEC0EAA5560044808AA6BB002EF6EE807BEFF6E5B3EAAA";
    attribute INIT_37 of inst : label is "C34E22F60F4768FE278DAC303410046BABB07087D749D125560FAEDBBF05FAED";
    attribute INIT_38 of inst : label is "A1F05AA8F4F0FABE0BC26AE0E209F447DB4AD31D131EDAEB48EA8BBED2348C34";
    attribute INIT_39 of inst : label is "9B82BFE9EBDAFFBCA666EE222A6D2D2ECAA55CB2D2E2AC2F8A88563C23D3882E";
    attribute INIT_3A of inst : label is "F83EA0BBFB0BBF6FD42EFDBF50BBF6FD02EFDBF40BBF6FD02EFD500BBF6E6F9A";
    attribute INIT_3B of inst : label is "7A1A86D6967CAA182A86299F99D86A57CD3E22138F078577D0FA9BBFB0AF769A";
    attribute INIT_3C of inst : label is "20EF8BE072F818BE0ED45478D51354DF5D785844BE2A621B0AA525E5A18167D6";
    attribute INIT_3D of inst : label is "C12701E8F130ED1E701D30EDC0BC303EF8BE0F2C308A8E8F8FE232F018BC0BC0";
    attribute INIT_3E of inst : label is "30EBCC209EA0C2F30C209C6ACB0BF08301AB0CB08030C209C6ACB01AB0CB0809";
    attribute INIT_3F of inst : label is "B0A7BF0C207A3C1AB2C308846ACB0C207A3C1AB2C30881AB2C30864FACB0C9C0";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "9D5AC5B546DB6263DF85C4B48F92D23E555500000000000000008A6770F1FBE2";
    attribute INIT_01 of inst : label is "0D6794CBF1E7163C21C3271EB899DCB89BC12004A455EFE7E3FDD59193C77C17";
    attribute INIT_02 of inst : label is "E6C6950000783300441010406AF22029AAF1AC6BDEC7BD1AF1AEFFE49207BC78";
    attribute INIT_03 of inst : label is "9E36778D9DEBC6372B7E6B359C8CBECD6FCB1A00CF04C9CB525632F9C5BFEB3E";
    attribute INIT_04 of inst : label is "C521555A34A71675A5995C564EA0FC2484984BD96C925F1FAEC2C1D9EF76BADD";
    attribute INIT_05 of inst : label is "976A41260176A92D59A96477966A81F671AC5D8A8E75F1DA39D55A878054ABD9";
    attribute INIT_06 of inst : label is "E5A595F7105AD586764554ABAF9A81DB1002ADD4C9D75B52ADD59AA0FC59AA4C";
    attribute INIT_07 of inst : label is "4B4A890706A25540A9BA5E9FA5E93A4E8964778AA80A42932545C6F699555555";
    attribute INIT_08 of inst : label is "5655A83F15A6D552A0510FC2AA814C8A84C9D72A1325568145322A6CA9BA2051";
    attribute INIT_09 of inst : label is "3BD7E74C0E0290245A1E87B3B2FB771881F1F3932325FBE72C2CE6844285D151";
    attribute INIT_0A of inst : label is "C6F7EFCBE46BD4EDD6BB9C0BC0FBE76FBDDAEB667BD9CEF76FBF9B47F32FBE67";
    attribute INIT_0B of inst : label is "F770737BBE0805773EDD9DBAF767BCA35DF3DD9EC28D756FBE0B467D19F44BFE";
    attribute INIT_0C of inst : label is "FB5FB769894218561D9D6875E77E3E75FD783EDD37AD30CDBDB0C1FFF410FFC6";
    attribute INIT_0D of inst : label is "82D0C9732F8C9CBCBEF9DCD1DDBDD9EF7677D9DE3677ADDAEB7675F14D49683C";
    attribute INIT_0E of inst : label is "3E102FCF8C0BE33EF9D5EF44B8EE8B30D3A1D8EF76B7F17DFBB6C93E801F0C9F";
    attribute INIT_0F of inst : label is "BBBBBBBBB9B999999999BBBBBBDFE8387EED7EEF3F65752E38B45413CF4B8E7A";
    attribute INIT_10 of inst : label is "999999999BBBBBBBBBBBBBB9B999999999BBBBBBBBBBBBBB9B999999999BBBBB";
    attribute INIT_11 of inst : label is "8511BBBBBBBB9B999999999BBBBBBBBBBBBBB9B999999999BBBBBBBBBBBBBB9B";
    attribute INIT_12 of inst : label is "EC834B4BF3F4C35CCCEC8FF88C6D239D34855FC631DDAFE6D9524F3FFB540F4B";
    attribute INIT_13 of inst : label is "14F55FFDF1C5232A799BC6DEA99FBCF1F8D65DB33021212393955FF3B23157FF";
    attribute INIT_14 of inst : label is "3396786B86F963A67A6B96F863B67A7075C41DB932C7B954ACC47971E655A833";
    attribute INIT_15 of inst : label is "F378DCFCDFE58816685FC03950E9702CCFCDC090E1B97331C0384C0BFCEEB300";
    attribute INIT_16 of inst : label is "F96011CEC0BCF3370243E5C862D00BF2F75BFF3B3330263DE6CDEE32E2C40B07";
    attribute INIT_17 of inst : label is "6A9BF0C495CF3E58060C0B3F37E58150E5302CCFCDC09F96021F3E58053C0B3C";
    attribute INIT_18 of inst : label is "B0301601EB034B438B8CFC47F193C44F197C45F19F31FF3A7E8C4B2025FC833E";
    attribute INIT_19 of inst : label is "50D5B08F842BB129D99604B0F92CABCCF1ED65B70FC9FF741A01601ECCB741A4";
    attribute INIT_1A of inst : label is "59DE376BCEF7C45276FCD5F7967FEDD8FB599697921E31F1A620329BAF1D530A";
    attribute INIT_1B of inst : label is "0CD0D35B0B970F251ACC69A59FF561D55555D556296902C49680B3F5C132C1EF";
    attribute INIT_1C of inst : label is "61AC6BDB8856A92F7E557C1F9197B98F37FFD59AF9197BBDFC1F9197B9F34687";
    attribute INIT_1D of inst : label is "49E706FC0A7B67755659BB128DDAFE730998E7C56C7B30DCC56DB87F9126579F";
    attribute INIT_1E of inst : label is "8E0297C18F0255F3644A3B8CD912778EE2FDD127C9E3D5645E65FACE1E767B9C";
    attribute INIT_1F of inst : label is "D56CDD4DDB355AD3543BD50CF543BD50CC611EF712F96CD156C565B456595BC4";
    attribute INIT_20 of inst : label is "3838383A7BA838F8F8787870F8B8B8B93A7AFAFABB3B7F9A5B2C7CD56FFFF1AC";
    attribute INIT_21 of inst : label is "4454554C54555454471A6C649AB940531D7C915515551110D79F245545D10428";
    attribute INIT_22 of inst : label is "A6F6498B5405D561451565551565551565551561C69B1D347AF40F54450C5455";
    attribute INIT_23 of inst : label is "766FE6E954E54454454455455455855455555C50C54C54C5455445505505507D";
    attribute INIT_24 of inst : label is "5561571571571B69ADD37285034981DA7F79FFE59407FE68E6CDA7DE721A48FF";
    attribute INIT_25 of inst : label is "961A68649AA94406B55045544956157157157155154155151551144154154157";
    attribute INIT_26 of inst : label is "5465465475465151551D51151551D55555555955555555954554554954554554";
    attribute INIT_27 of inst : label is "DE0A1B95C07FFE4FCC696924925C5567FDD54544446557557556557557546547";
    attribute INIT_28 of inst : label is "259E49669EF3205C0C84921A49D5FF741B1E3FFE7E7811BCB64E937FFDBDFFF6";
    attribute INIT_29 of inst : label is "74B77EF5C21DB305B0D83580DD2FBD3306C360D60374BCBDB3075B0D6037FF69";
    attribute INIT_2A of inst : label is "D60E09F6CC47234CC00CD2F4C36CC16C360D60374AB5AAC360DFF36CC1B0D603";
    attribute INIT_2B of inst : label is "C288C883D574D6CDB03ABC0DB771C15230C8DB3012F4BABF595ACB5DC89F6CC4";
    attribute INIT_2C of inst : label is "CDB30148A7ECC012EFB12F125552330322111033FFB9733212220F3311443513";
    attribute INIT_2D of inst : label is "E77DF7ADF4F01FFF93F31AFDF626E26AE36EAEEF6CC07FFFB012883CF3F1F2F3";
    attribute INIT_2E of inst : label is "429AA83F0EB6EA10F0F73099B8967ED453191DC2AD0128BA80D74465642BD36F";
    attribute INIT_2F of inst : label is "678D549D7767ADDBEF7638D1445E767ADDAE32B945098B653F6E880BF3081B8A";
    attribute INIT_30 of inst : label is "BEE6FCD4AC4CBE09E0223110C2252D30232FBCD4AC524E6C0B03193D2B1DAE37";
    attribute INIT_31 of inst : label is "BE065701BD1F0AF4A30A4B4B2C4BA193C9CBED7E1865701B9B2E18CBE3A2F1AC";
    attribute INIT_32 of inst : label is "EE029D5CACFCF4A30A434B1CFB54BD6FD9DEB6778D55965567EE6CB86FA2F1AC";
    attribute INIT_33 of inst : label is "AEE88F42AEA00F0EB6EE88F41D7E97D730BFF44A58ACB04A687BFF7425837B8D";
    attribute INIT_34 of inst : label is "36E7F7DF9DDF4E7FF3AC0FCB4C6BCB4C6BCB486BCB4862CE06D5FA70FF7CDAAA";
    attribute INIT_35 of inst : label is "5A33D54581ACCF7411D66B1770CFF965AEF3B59C26F7560AFD9DDBE699455909";
    attribute INIT_36 of inst : label is "05A5916435A257469188689F5554A9552A2C555DAA9827586A675FFBF3D76AA8";
    attribute INIT_37 of inst : label is "59B5B16791006117ED94F8A2648B220A8FDB123FDD9BF9BA55AA75156EA5A7B1";
    attribute INIT_38 of inst : label is "B5673D075A8D10071D9DF44C49C35AF17E386B16A616AD61FC7331045A1E86AF";
    attribute INIT_39 of inst : label is "1568165191551A361515511DD59F76E5B00C9FD5766273C90B877119DD7D6C87";
    attribute INIT_3A of inst : label is "9E9B4AD16EA56E591A95B9646A56E591E95B9647A56E591A95B9F6A56E57515C";
    attribute INIT_3B of inst : label is "1F17C311680B3E134FC4F0440C5E20D4F7D5B2F1216565555A6D1D16EA445415";
    attribute INIT_3C of inst : label is "35498263967FEDD8F3D6DEBC05801EFFF756EE6D95B76F10F831E121E17F1133";
    attribute INIT_3D of inst : label is "7BF1ED5B0AED4AD61EC66C6A48C49AD49C2611479A87C732327BD6778D149DBF";
    attribute INIT_3E of inst : label is "5A43868C35FC78E1A6AC37776D739AC1ADDDB7DE8B1A6AC37776DFDDDB5DECBC";
    attribute INIT_3F of inst : label is "174559E7B355C2DDDB7DECFF776D77A355C2DDDB5DE8FDDDB7DEC70544DF7C7A";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "E9CFCEC186D20000C8BF0EAECAF2B32B11005555555555555555408D6989AAA0";
    attribute INIT_01 of inst : label is "6FEF9BA9CFF63FAD92DABB337361054042A7319ECF4052AEA0011CAD180CC8B0";
    attribute INIT_02 of inst : label is "1586C088008C0B0804F4ECEF8DFC24E227CF6ADDF6ADEEF6AB7502AEB27DAADC";
    attribute INIT_03 of inst : label is "B28664819B286600926A68DDB88D6B28F188FE702DFC25B276F625AFCDD00EAB";
    attribute INIT_04 of inst : label is "B2C6AAA56862C9A7D890A8309B4DA21B1A698606006C669C19AB09DA2074491D";
    attribute INIT_05 of inst : label is "28BD0C22D2ABD168A2F528622ABD0DA0ACA0A2C5782880CDE0AAA5061C185628";
    attribute INIT_06 of inst : label is "40DC8E6C1A65988A28B3A854888575881B4959C9864E867159CA2F4DA2AAF4B1";
    attribute INIT_07 of inst : label is "5A25465A7151AA9656A5996A5B96E599452862255695B56C489682A168EAAAAA";
    attribute INIT_08 of inst : label is "E22AD368A8028AA15432DA2955DEB1057B124E1DEC4AA950CAC4958056851432";
    attribute INIT_09 of inst : label is "0200097CCBBBCEFB1CC7B0CFA1ACD68A8A08BF225359AEAFB088D1775178B1F1";
    attribute INIT_0A of inst : label is "64000086BC60A581D0C201A216AEA76801D80064011980876431DC410A1AAB66";
    attribute INIT_0B of inst : label is "41AF4E420127302800257900074C3AC41D161D30DB10740020F814E0528178A0";
    attribute INIT_0C of inst : label is "02400959B54FDD7A0753A374CCBC437459E20025A4824529A2C721A2821D2864";
    attribute INIT_0D of inst : label is "82AC2E331ACD5D6C6BAB5A3100C1DB08760819920664A1D12476C819A00BF8E3";
    attribute INIT_0E of inst : label is "0BF5ABAAC996B2AAADD92474C1380E822AE1DA08744A19A00026E5FE30C9C2C7";
    attribute INIT_0F of inst : label is "222222222023333033333222324A201B40092D39604482ECD442D68624BA316E";
    attribute INIT_10 of inst : label is "3333033333222322222222202333303333322232222222220233330333332223";
    attribute INIT_11 of inst : label is "B048222222220233330333332223222222222023333033333222322222222202";
    attribute INIT_12 of inst : label is "8A18787ED0A09DD8AACA02A8BA71EEBAA5800466C85DB077157E042068D698BA";
    attribute INIT_13 of inst : label is "8784040109B561BDF11BB717F74F248DA81155C2ED1571FE9EC4040A28190103";
    attribute INIT_14 of inst : label is "C6472676E72472776E72476C76C725474107D1E12B8461A04BAA61A11C6811EA";
    attribute INIT_15 of inst : label is "6C16441ACC1DAA43BB6B067446DDE374B1A28DC6F9F4512EBDBC78DD00F93CFB";
    attribute INIT_16 of inst : label is "C76BC8C68DDA12C3371B1DA30AC8DD00914442832CB3716555C4D3CF4EC3DDF0";
    attribute INIT_17 of inst : label is "2D57CCBD1046B1DAF298DD068B1DA446D12374B1A28DCC76BC86B1DAF2B8DD1A";
    attribute INIT_18 of inst : label is "EEE59B19BBAB2FAF2BA42BF7AFD6BE6AF96BF6AFDA9914F59E6E7F5E25405101";
    attribute INIT_19 of inst : label is "5B354D823F763413172F68DCFAB6110343B77DF1033D9FC59B59B19B4BBC59BF";
    attribute INIT_1A of inst : label is "5992074010C43C73760819B5D66CA1D928EBE7DDBE383B8062DA82DFEE9354DD";
    attribute INIT_1B of inst : label is "F4EECFEA97E550969A236F6EC00455000400C4008E7D3B3CDA3D9F6CD0ADC77B";
    attribute INIT_1C of inst : label is "636ADC56261413AB58101F105D40756601001EB705D404310F105D4075E43673";
    attribute INIT_1D of inst : label is "EFA83B63DC8A66467A9E033F81D64D44DD9200C7AFC8F1DC01414319E3F46C22";
    attribute INIT_1E of inst : label is "CAF7348EECF7A44B6CFE43801B3F2C80EE01F3F1C90017BC7F64801AF77403B0";
    attribute INIT_1F of inst : label is "2942E9425705EF85AD6C6B5A1AD646B58372B7B63FABA21A7AF3BE877A9CECCE";
    attribute INIT_20 of inst : label is "89A9A98A68E949EB2BEB6B6BE3EBEBE968EAAAAA882AA210ECAAC017B8AAAD1D";
    attribute INIT_21 of inst : label is "5CF5BF5CF5BF5CF58F3CFCDF75FBE1FFFDFEBF5FF5FBBDDBCF3F2DD7EFDBF669";
    attribute INIT_22 of inst : label is "CF5DF75DFE16FD77F63D7FD73D7FD63D7FDF3D737D35FFFCF554DFF59FDCF7BF";
    attribute INIT_23 of inst : label is "AA685A0E83EF7BF7FF7FF5FF5BF5FF5BFFEF59FFDF7DF7CFFEF79F59F59F58D7";
    attribute INIT_24 of inst : label is "BD77DD7DD7DD3ED37BFFF5D70DDB25786CE1A129846D82AF6A3F847B28FB46D2";
    attribute INIT_25 of inst : label is "DF3CFCDF76FB6F1FAFF5F5FE6BD7FD7FD7FDFFDFFDCFDFFFFBDE7F67D67D63F7";
    attribute INIT_26 of inst : label is "7FE7F77F67F671F7DF79F51F5DF59FFDFF9FFDFDDFD9FDDFFDFF9FFDFDDFD9FD";
    attribute INIT_27 of inst : label is "3806940013B7FF3D0F59DBCF35FDFFCF7FFDFDC6B9E7DF7DE7D67D77D67FF7FE";
    attribute INIT_28 of inst : label is "8808B24B2C5681B00A52D8C079C079B8D4709022E2E03909A23BAE68A149A285";
    attribute INIT_29 of inst : label is "4A0340864CC546800291A41A92820546800A46906A4A0A254683402906A44032";
    attribute INIT_2A of inst : label is "566C2D151A008D51A00AE802F151A001A42906A4A00A200A4690FD51A002906A";
    attribute INIT_2B of inst : label is "070CBD08002768A504089A414368831F687250681F0A018E595CA2CD42D151A0";
    attribute INIT_2C of inst : label is "F50680320181A0560C23773F00088B89B99B9989020E76AAAA8AAE6AAB223489";
    attribute INIT_2D of inst : label is "F4630BE10C11B4AA9A1683A048D861415A56000941A010088E1C23F000CEDC63";
    attribute INIT_2E of inst : label is "AFB998C33FF782EB8C164FDBBFD5509E69FC11CFF101F8E0BC3CA3C547EF14D1";
    attribute INIT_2F of inst : label is "68731A23C74491D21076C439EC7F75091DB1CC9DE7A5FC7917780CB464FC5EB5";
    attribute INIT_30 of inst : label is "6B65F35734786BEBCFB32F4F3B97EDCBBE1AF357347EE663E8F0EADDEADDB147";
    attribute INIT_31 of inst : label is "6B3A53BEC8C33B77A0BBE2F8F8FF4EAFD7D6A56BCBA53BED98E9FE96B7BEADD9";
    attribute INIT_32 of inst : label is "0AFBA007234C77A0BBE2F8E8A95FD3A019928664819EA703B38663A7FFBEADD9";
    attribute INIT_33 of inst : label is "1380F808396CB8FFF5380F80856A19128FD44C7BEB63B3F7F80C40E73EAC8232";
    attribute INIT_34 of inst : label is "4D1C763072D0C1C40F8CCC2B0B742B03742B0B742B027C3E0F00565881580000";
    attribute INIT_35 of inst : label is "EAD631AE8FE358E7F17AF8C1A4274D540160C433D7077ABB01992077DE4051F9";
    attribute INIT_36 of inst : label is "EA5A00A16A5CC6754983778A3AA85599159A385B57490A08D5A13902160E7002";
    attribute INIT_37 of inst : label is "E94E8F023D194BDE09849A28C357D5512A3404E1FFCF43D6F55220A8285A220A";
    attribute INIT_38 of inst : label is "8D4063845B93AED4DD038768FFC75A0562426AC6DCB04449866CB5D468DABE8C";
    attribute INIT_39 of inst : label is "E994DC3A2CE3906DD59D5D59197475D7C55A4752444FC125BB3B2B923D63AF76";
    attribute INIT_3A of inst : label is "B970E5B1285828A82960A2A085828A82960A2A085828A82960A20458288E8469";
    attribute INIT_3B of inst : label is "D19B22F478F8B09A5C26A6B46B783813861E8EF3F273B11005C3AB1285B58A60";
    attribute INIT_3C of inst : label is "0665B94DD66C11D10C0F0FB8D3930E40047A38411ECC1E904E218D2D29AEAD2A";
    attribute INIT_3D of inst : label is "FECF7354DDCC14BEF7C58D14C82CF6A65396F9EDBEB333A5A5DED664831CDD82";
    attribute INIT_3E of inst : label is "9F4D8DCC75D8EF637D887660D30CBEB3F9834E3EB637D887660D389834C3E3F3";
    attribute INIT_3F of inst : label is "3CA0C3ED8CD4379834E3E3B260D30FACD4379834C3EBB9834E3E30C1BE30F3DF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "AEEADEB9A6DFBBBBAF0FCE9EBBBA7AEE44440000000000000000869A7F299AE0";
    attribute INIT_01 of inst : label is "DBEEAEC3F3AB7EB36EF7EB7E2A6E367B00DFAF7E8A4442EAE1144EBA1DFEBF6D";
    attribute INIT_02 of inst : label is "D7DE93BBBBE296BBBF8F8FAAE304DE5F8CBBA9E8BA9E8ABA27A4126EBA2E89EB";
    attribute INIT_03 of inst : label is "FF2B7BEADEFAE767C86EEB9EAB876EE6EDBBBAEBD42FEDE87ABA1DBBDE91C66E";
    attribute INIT_04 of inst : label is "FEFFAAA5FA7FF9BF5FFFEFFFBD7FFF9BFE6FA7E6FE71ABA9CBECFEDCF2B77FAD";
    attribute INIT_05 of inst : label is "EAA5FFFFFEAA5FFFAA97FBFFEAA5FFFFBFFFAAA56FFBFFF5BFEAA5FFFFFE57EF";
    attribute INIT_06 of inst : label is "FF5FFEFFFFF5FFFBFBFFAA56AAA57FFFFFF95FFBE6FFA7F95FFAA97FFFAA97FF";
    attribute INIT_07 of inst : label is "FFE566FBF959AABE56E5B96E5B96E5B967FBFFE557F5BD7FFBFEFFFD7FEAAAAA";
    attribute INIT_08 of inst : label is "EFEA5FFFEFFFFEA95FFEFFF955BEFFE56FFEFF95BFFAA97FFBFF95AE56B59FFE";
    attribute INIT_09 of inst : label is "BF935C4F3DCE739CC739CE7239B9A6DE8CFFF2FBD79ABA6ACFFDBD7FFD6FFFFF";
    attribute INIT_0A of inst : label is "E72754E6E873E5B6D76EDBFEF99A6B7BCADCFAB73FADEFEB77EA99451399AEB7";
    attribute INIT_0B of inst : label is "257097D2C985B17F35711ECF4B76F1F22D23ADDBF7C8B536EFBBC6FF1BFC7AFC";
    attribute INIT_0C of inst : label is "A85D5C6DEB7A197A1613EEB4B6F327B44F2D3571F4CFE8FDCFE8F9FFF392FFE7";
    attribute INIT_0D of inst : label is "A3F3DA6F9BAF7E6E6E9A9B61CD86DCFEB73FADEFAB7BEADDFEB7FFB9E92AF8EF";
    attribute INIT_0E of inst : label is "3FBC7EDBB536EC26BADDBBB77C8BAABDBEA2DCFEB7FFB9E9D584AD8AEABC3CA6";
    attribute INIT_0F of inst : label is "FFFFFFFFFEFFFFFEFFFFEFFFEFBFFBFBF5617D5A3987E7BBA73F87D1BBEFE9EA";
    attribute INIT_10 of inst : label is "FFFFEFFFFEFFFEFFFFFFFFFEFFFFFEFFFFEFFFEFFFFFFFFFEFFFFFEFFFFEFFFE";
    attribute INIT_11 of inst : label is "E4FDFFFFFFFFEFFFFFEFFFFEFFFEFFFFFFFFFEFFFFFEFFFFEFFFEFFFFFFFFFEF";
    attribute INIT_12 of inst : label is "BEFBF9FAC179F2DF99BEE098FFEFEE8A6F8545E7FD6DDCA65B7A0561B687C6EE";
    attribute INIT_13 of inst : label is "D3B11514F8E3E3422CC6EECC0AECF3F09846DFBF7BDBEBEEAE911452FBB15114";
    attribute INIT_14 of inst : label is "BFC7BC7BC7FF7FC7FD7BD7BD7BC7FF6F14E3846CA6E038FF02EF6CB80E3FC3BA";
    attribute INIT_15 of inst : label is "BE0F141DBC75FE930CAC3DBC4D71F7E56153DF8D71DF514BF35D7DF9458BF3BF";
    attribute INIT_16 of inst : label is "4D7BBC5ADF99158F7E3535AA3FFDF951CC9D574E68F7E2733EDBFC3B3FDFF8E4";
    attribute INIT_17 of inst : label is "02EF1BDB6146535EE3FDF9074F35E88D71B7E52193DF84D7BBC6535EE3CDF915";
    attribute INIT_18 of inst : label is "3B0F7AF7AEEEEEEEEAE4FAF7FBDFAF6FBDBAE7FB9471F425F44FFD7FC751B113";
    attribute INIT_19 of inst : label is "DFE7BF8FCBE39FC2D3BCCE35B38CC15E53430C454FE22FC77AF7AF7A5AFC77AD";
    attribute INIT_1A of inst : label is "6DEFAB7BEBFEC87EB73DA1D69B7BDADDF2FA865FBA0BBFB0BED8BBBA8B9E7FFA";
    attribute INIT_1B of inst : label is "CBF3F2FA768608B73EDDFBEF811A5D9111129112986525CFB8CFA22FA7FDDBAD";
    attribute INIT_1C of inst : label is "A3A9EB53A69EC3ED69444B956D556DCAB5114FBE56D562E9AB956D556DAF78CF";
    attribute INIT_1D of inst : label is "FBF27EFCFB7FB7B87EEB2F7AEAD76B73FADDB7B7EEFB961561FBFF6E97A87ADF";
    attribute INIT_1E of inst : label is "AF3E87DFBB3EB7BFB5EBEFF92D7A3BEBF3A2D7A3DFB7C7F97EB7ACFF3EB7EFC9";
    attribute INIT_1F of inst : label is "2DFFADFE5F71FE8AB3AFACEBEB3AFACEBF57FAD57A9BE25A7EE3EF887EE8FADF";
    attribute INIT_20 of inst : label is "3E3E3E3EFEFEFEFE7E7EBEBE3EBEBEBE7E7E3E3E7EBE7E65FF1EFDC7FFFEFD7A";
    attribute INIT_21 of inst : label is "AAAA2AAAAA2AAAAA26E5BB9AAAACAA6A26B8DAEBAEBAAAAAA96EB6BAEAAAAABE";
    attribute INIT_22 of inst : label is "5B99AA8A8AABAAAAABAABAAAAAAAABAAAAABAAA9896E262AAA82AAAA2AAAAA2A";
    attribute INIT_23 of inst : label is "B699BA6AA6EAA2AA6AA2AA6AAEAAAAAEAAEAAEAAEAAEAAEAA6AA2AA6AA6AA666";
    attribute INIT_24 of inst : label is "AABAA8AA8AA89B96EE62A292A9FAD97A76E9F92DA79AFADCADCBB5FB7FFB79E5";
    attribute INIT_25 of inst : label is "A665B99AA8A4AAA6C6BAAAAA9AABAA8AAAAA9AA9AABAA9AA9AA8AA9AA9AA9AA8";
    attribute INIT_26 of inst : label is "AABAA8AA9AABAEAA2AA6AAEAA2AA6AA6AAEAAAAA6AAEAAAAA6AAEAAAAA6AAEAA";
    attribute INIT_27 of inst : label is "CB82FF1451386CCAAEA9625B6EE6BADBA22AAAAAAAAAABAA8AAAAABAA8AA8AA9";
    attribute INIT_28 of inst : label is "59698659656B9EBFF5A21B9FEA914AB5BB0BD16EAE2E3FBBAEEBB87BBBF1EEAF";
    attribute INIT_29 of inst : label is "5A494B9FFF9BFBB1CE5F94E65692EBBBB7397E53995A4EEBFBB95CE539955196";
    attribute INIT_2A of inst : label is "BA9AA12FEE34BAEEEFF5A90BC2FEEC7397E53995A6896E697A56CAFEEDCE5399";
    attribute INIT_2B of inst : label is "0EBADA7A850C65EBBBCBAEB3F97C7E3ABBBFBBBBFA5A4B97EAEBEEE5BA12FEE3";
    attribute INIT_2C of inst : label is "2BBBBD6FF6BEEFFA38F7AF7A113BBBAABAABBAB916E86E6F77776AE6F6DDEB31";
    attribute INIT_2D of inst : label is "AFEB7ABFADDE6839B22B8AFD4E9B59EC5956E3BAEEEF111BBA5BEEF553BBCBFE";
    attribute INIT_2E of inst : label is "FFAAA8F97EA4AEBFAEE3AFCAFCBE521B4DFDAFDFA52DF82BAEBFF3F7E7FAFEEF";
    attribute INIT_2F of inst : label is "7BAA9FEFEB77FADCEEB7FBAD397EB6AFEDDEAFA9B6EDE961184AEBFABAFE12AB";
    attribute INIT_30 of inst : label is "6EA59CA7EB7E6EFA73EAF6DEFEB7BFB7EB9B9CA7EB7EBA6EFBBEFAA1FAADCEEB";
    attribute INIT_31 of inst : label is "6EBEAECF9EFD7E87EF3EBAFB8DFADFABE7F66A6EFBEAECFA9BBE28E6EEABF2BF";
    attribute INIT_32 of inst : label is "FF3EED47EE7D87EF3EBAFB8D9A9F93E06DEFAB7BEA1FBA43E21A6EF8AEABF2BF";
    attribute INIT_33 of inst : label is "B0BABA3ECAEBEF3EA64BABB7DA66AA47EFFF487EFBEEECBEF83B4597EFBB3FCC";
    attribute INIT_34 of inst : label is "FEEEEEF7AABBDE641FBDB8EF3C28EF3C28EF3C28EF3C2EBE8FD061FC922F8AAA";
    attribute INIT_35 of inst : label is "FBB1E9FFBBEEC797A1BEFB856FD90BE4F5BF85FFE7FB7EEDC6DEF2A65844FDFF";
    attribute INIT_36 of inst : label is "FA5AFFBFFA5BFFFD7FFFD6FFFAAA56AA959FFBFE557FFBFF95BFFD4271D96AAF";
    attribute INIT_37 of inst : label is "FFFFBB52E9A67E9FE1A5AAEBEC46112CFFBB945B4F26EEBAA15FFFEFFF5AFFFE";
    attribute INIT_38 of inst : label is "F8731ACC7AEEDBE7ADCE686DEAD87A21EB3FEA8E8EBF0D7FBE7FE1E4EABAEFF7";
    attribute INIT_39 of inst : label is "EFD7FFFEFFEFFFF96AAEAEAAEA24B5B67FF1469A487BADEDEEEF061CFDEFEEA6";
    attribute INIT_3A of inst : label is "FD7FF5FFFF5FFFBFE97FFEFFA5FFFBFE97FFEFFA5FFFBFE97FFEAA5FFFBFBFEF";
    attribute INIT_3B of inst : label is "8F8EEF6D833BAF8FABE3CDE3DE0BBC47BECFBBE7AFA3E44445FFEFFFF5FFBBEF";
    attribute INIT_3C of inst : label is "686DAB6A9B7BFADDFEF030236C3DF044513E1B361FBA7F037F3878F8F8F078C7";
    attribute INIT_3D of inst : label is "FAF3EE7BF8A6F0F73EB4E7F0FBCFBEE6DEB7ADBFBEEEE2F9FDEB5B7BEA1FADCF";
    attribute INIT_3E of inst : label is "19485FBD878DEA17EFBD847FFBB97EE7E1FFFEBEE77EFBD847FFBB1FFFEBEEFC";
    attribute INIT_3F of inst : label is "3FF5D7EFBB9EFE1FFEEFEEB07FFBBFBB9EFE1FFEEFEEB1FFEEFEE321FEBBBCFA";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
