-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "B2AC7F73A0E0679BD9CABCC59633AFBED916B61BD2AD1FBEDFA029F6D44AE9E9";
    attribute INIT_01 of inst : label is "AD08988A366ADA35AD1B34B0DDAB6AA4DD9B42FEAB698FFFCF801ABEDD4765AD";
    attribute INIT_02 of inst : label is "2366C61B356B4CD451B834A8DC1AB70DC5AB5026A3706AD0A8D6B46E0D8C3706";
    attribute INIT_03 of inst : label is "DBE0A1425334A807DE8B82E44F525642F21798BD0DB72C94929261FFA2A376AD";
    attribute INIT_04 of inst : label is "5DA7E4BFCFC806E483725DB3393141C116AAF534F876290996CD54D8BA6B2482";
    attribute INIT_05 of inst : label is "BC8F3769B9FFFFFFFFF9361C4CD30991864D1CD4C322384A5010AE91F92FF372";
    attribute INIT_06 of inst : label is "7116D869AEF11E272FA1DBD299DA59B639FE4A45EE5BBEC4447895FE243252EC";
    attribute INIT_07 of inst : label is "4597367DF5FCFC25F997265C895224DBD36E47AD1EBD7BFBBFAFFF3E1054FCC0";
    attribute INIT_08 of inst : label is "C1A1842D00D8635B16861034376580056DB57589FDFDB18CDAF2CFF699A54D6D";
    attribute INIT_09 of inst : label is "55555555555555555555555578742E5534EE676CE79EFFFFFBCF386220B418C6";
    attribute INIT_0A of inst : label is "29BB4F3CF7FE926471987E788ED3FFFFD5555555455D55555554755555555157";
    attribute INIT_0B of inst : label is "F42E540CCFF429FE807E1F97B2E65C8A4CBEE0B47DC59205E45892445E44CBF7";
    attribute INIT_0C of inst : label is "AFB1D9B29CF7E2548616009A57CD73914EBC429AD12DF2837AA42265F3D416E7";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC11151200B27321FB1C022EBD929AE";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "B2AC7F73A0E0679BD9CABCC59633AFBED916B61BD2AD1FBEDFA029F6D44AE9E9";
    attribute INIT_11 of inst : label is "AD08988A366ADA35AD1B34B0DDAB6AA4DD9B42FEAB698FFFCF801ABEDD4765AD";
    attribute INIT_12 of inst : label is "2366C61B356B4CD451B834A8DC1AB70DC5AB5026A3706AD0A8D6B46E0D8C3706";
    attribute INIT_13 of inst : label is "DBE0A1425334A807DE8B82E44F525642F21798BD0DB72C94929261FFA2A376AD";
    attribute INIT_14 of inst : label is "5DA7E4BFCFC806E483725DB3393141C116AAF534F876290996CD54D8BA6B2482";
    attribute INIT_15 of inst : label is "BC8F3769B9FFFFFFFFF9361C4CD30991864D1CD4C322384A5010AE91F92FF372";
    attribute INIT_16 of inst : label is "7116D869AEF11E272FA1DBD299DA59B639FE4A45EE5BBEC4447895FE243252EC";
    attribute INIT_17 of inst : label is "4597367DF5FCFC25F997265C895224DBD36E47AD1EBD7BFBBFAFFF3E1054FCC0";
    attribute INIT_18 of inst : label is "C1A1842D00D8635B16861034376580056DB57589FDFDB18CDAF2CFF699A54D6D";
    attribute INIT_19 of inst : label is "55555555555555555555555578742E5534EE676CE79EFFFFFBCF386220B418C6";
    attribute INIT_1A of inst : label is "29BB4F3CF7FE926471987E788ED3FFFFD5555555455D55555554755555555157";
    attribute INIT_1B of inst : label is "F42E540CCFF429FE807E1F97B2E65C8A4CBEE0B47DC59205E45892445E44CBF7";
    attribute INIT_1C of inst : label is "AFB1D9B29CF7E2548616009A57CD73914EBC429AD12DF2837AA42265F3D416E7";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC11151200B27321FB1C022EBD929AE";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "B2AC7F73A0E0679BD9CABCC59633AFBED916B61BD2AD1FBEDFA029F6D44AE9E9";
    attribute INIT_21 of inst : label is "AD08988A366ADA35AD1B34B0DDAB6AA4DD9B42FEAB698FFFCF801ABEDD4765AD";
    attribute INIT_22 of inst : label is "2366C61B356B4CD451B834A8DC1AB70DC5AB5026A3706AD0A8D6B46E0D8C3706";
    attribute INIT_23 of inst : label is "DBE0A1425334A807DE8B82E44F525642F21798BD0DB72C94929261FFA2A376AD";
    attribute INIT_24 of inst : label is "5DA7E4BFCFC806E483725DB3393141C116AAF534F876290996CD54D8BA6B2482";
    attribute INIT_25 of inst : label is "BC8F3769B9FFFFFFFFF9361C4CD30991864D1CD4C322384A5010AE91F92FF372";
    attribute INIT_26 of inst : label is "7116D869AEF11E272FA1DBD299DA59B639FE4A45EE5BBEC4447895FE243252EC";
    attribute INIT_27 of inst : label is "4597367DF5FCFC25F997265C895224DBD36E47AD1EBD7BFBBFAFFF3E1054FCC0";
    attribute INIT_28 of inst : label is "C1A1842D00D8635B16861034376580056DB57589FDFDB18CDAF2CFF699A54D6D";
    attribute INIT_29 of inst : label is "55555555555555555555555578742E5534EE676CE79EFFFFFBCF386220B418C6";
    attribute INIT_2A of inst : label is "29BB4F3CF7FE926471987E788ED3FFFFD5555555455D55555554755555555157";
    attribute INIT_2B of inst : label is "F42E540CCFF429FE807E1F97B2E65C8A4CBEE0B47DC59205E45892445E44CBF7";
    attribute INIT_2C of inst : label is "AFB1D9B29CF7E2548616009A57CD73914EBC429AD12DF2837AA42265F3D416E7";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC11151200B27321FB1C022EBD929AE";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "B2AC7F73A0E0679BD9CABCC59633AFBED916B61BD2AD1FBEDFA029F6D44AE9E9";
    attribute INIT_31 of inst : label is "AD08988A366ADA35AD1B34B0DDAB6AA4DD9B42FEAB698FFFCF801ABEDD4765AD";
    attribute INIT_32 of inst : label is "2366C61B356B4CD451B834A8DC1AB70DC5AB5026A3706AD0A8D6B46E0D8C3706";
    attribute INIT_33 of inst : label is "DBE0A1425334A807DE8B82E44F525642F21798BD0DB72C94929261FFA2A376AD";
    attribute INIT_34 of inst : label is "5DA7E4BFCFC806E483725DB3393141C116AAF534F876290996CD54D8BA6B2482";
    attribute INIT_35 of inst : label is "BC8F3769B9FFFFFFFFF9361C4CD30991864D1CD4C322384A5010AE91F92FF372";
    attribute INIT_36 of inst : label is "7116D869AEF11E272FA1DBD299DA59B639FE4A45EE5BBEC4447895FE243252EC";
    attribute INIT_37 of inst : label is "4597367DF5FCFC25F997265C895224DBD36E47AD1EBD7BFBBFAFFF3E1054FCC0";
    attribute INIT_38 of inst : label is "C1A1842D00D8635B16861034376580056DB57589FDFDB18CDAF2CFF699A54D6D";
    attribute INIT_39 of inst : label is "55555555555555555555555578742E5534EE676CE79EFFFFFBCF386220B418C6";
    attribute INIT_3A of inst : label is "29BB4F3CF7FE926471987E788ED3FFFFD5555555455D55555554755555555157";
    attribute INIT_3B of inst : label is "F42E540CCFF429FE807E1F97B2E65C8A4CBEE0B47DC59205E45892445E44CBF7";
    attribute INIT_3C of inst : label is "AFB1D9B29CF7E2548616009A57CD73914EBC429AD12DF2837AA42265F3D416E7";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC11151200B27321FB1C022EBD929AE";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "41B8EC4AA2AD486001D143C12AA4D844AACB2AE821D1A40B2038D61526A91036";
    attribute INIT_01 of inst : label is "36B2E45EBAF12E9D120D795EEBC4817B42440503FFB2AA1544889BCB2798AAF6";
    attribute INIT_02 of inst : label is "E0AD2BD569B75F6290DE797AEF3C49EEF3C4BFFBEABCD3617A74D8179A57ABCD";
    attribute INIT_03 of inst : label is "2DB9C2BC063166162C542507A2F1A9950DAA659276218A204408ACFD05EABD36";
    attribute INIT_04 of inst : label is "06082E08905DA82ED4971418EE3D14F153332C1A08A8D21A002A6A294AA8A8C7";
    attribute INIT_05 of inst : label is "45D08D6564FFFFFFFFFA10C48539108C4E2BC86A255D9800429485BA0B830497";
    attribute INIT_06 of inst : label is "82276792C9422AEA5B4014BCE47704D6E4FEDEE257E4874CE1FBB8FE4E031701";
    attribute INIT_07 of inst : label is "D6BC2436496B456CFA64C183264C19026080902601EB9080B800064D2C8B0D38";
    attribute INIT_08 of inst : label is "12D50B321164B46459542C5A4AAAE227B2BCBDAA6A36FA28032C225912E790B1";
    attribute INIT_09 of inst : label is "CE6666662746E6666662746F7F1678665620156D18BBFFE40412D0B446CB2D0B";
    attribute INIT_0A of inst : label is "628B297C012208198005818462CAFFFFE4BE61E334CE6666662666E4B0618532";
    attribute INIT_0B of inst : label is "0313E9F12009D0013B01A0BC1782F050810039BF0E6984668285606282E8104E";
    attribute INIT_0C of inst : label is "501A324CD7013426A6DEE764990E682091011419BBC4F128F04C0253E3140203";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4051400884880A236194C00021242";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "41B8EC4AA2AD486001D143C12AA4D844AACB2AE821D1A40B2038D61526A91036";
    attribute INIT_11 of inst : label is "36B2E45EBAF12E9D120D795EEBC4817B42440503FFB2AA1544889BCB2798AAF6";
    attribute INIT_12 of inst : label is "E0AD2BD569B75F6290DE797AEF3C49EEF3C4BFFBEABCD3617A74D8179A57ABCD";
    attribute INIT_13 of inst : label is "2DB9C2BC063166162C542507A2F1A9950DAA659276218A204408ACFD05EABD36";
    attribute INIT_14 of inst : label is "06082E08905DA82ED4971418EE3D14F153332C1A08A8D21A002A6A294AA8A8C7";
    attribute INIT_15 of inst : label is "45D08D6564FFFFFFFFFA10C48539108C4E2BC86A255D9800429485BA0B830497";
    attribute INIT_16 of inst : label is "82276792C9422AEA5B4014BCE47704D6E4FEDEE257E4874CE1FBB8FE4E031701";
    attribute INIT_17 of inst : label is "D6BC2436496B456CFA64C183264C19026080902601EB9080B800064D2C8B0D38";
    attribute INIT_18 of inst : label is "12D50B321164B46459542C5A4AAAE227B2BCBDAA6A36FA28032C225912E790B1";
    attribute INIT_19 of inst : label is "CE6666662746E6666662746F7F1678665620156D18BBFFE40412D0B446CB2D0B";
    attribute INIT_1A of inst : label is "628B297C012208198005818462CAFFFFE4BE61E334CE6666662666E4B0618532";
    attribute INIT_1B of inst : label is "0313E9F12009D0013B01A0BC1782F050810039BF0E6984668285606282E8104E";
    attribute INIT_1C of inst : label is "501A324CD7013426A6DEE764990E682091011419BBC4F128F04C0253E3140203";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4051400884880A236194C00021242";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "41B8EC4AA2AD486001D143C12AA4D844AACB2AE821D1A40B2038D61526A91036";
    attribute INIT_21 of inst : label is "36B2E45EBAF12E9D120D795EEBC4817B42440503FFB2AA1544889BCB2798AAF6";
    attribute INIT_22 of inst : label is "E0AD2BD569B75F6290DE797AEF3C49EEF3C4BFFBEABCD3617A74D8179A57ABCD";
    attribute INIT_23 of inst : label is "2DB9C2BC063166162C542507A2F1A9950DAA659276218A204408ACFD05EABD36";
    attribute INIT_24 of inst : label is "06082E08905DA82ED4971418EE3D14F153332C1A08A8D21A002A6A294AA8A8C7";
    attribute INIT_25 of inst : label is "45D08D6564FFFFFFFFFA10C48539108C4E2BC86A255D9800429485BA0B830497";
    attribute INIT_26 of inst : label is "82276792C9422AEA5B4014BCE47704D6E4FEDEE257E4874CE1FBB8FE4E031701";
    attribute INIT_27 of inst : label is "D6BC2436496B456CFA64C183264C19026080902601EB9080B800064D2C8B0D38";
    attribute INIT_28 of inst : label is "12D50B321164B46459542C5A4AAAE227B2BCBDAA6A36FA28032C225912E790B1";
    attribute INIT_29 of inst : label is "CE6666662746E6666662746F7F1678665620156D18BBFFE40412D0B446CB2D0B";
    attribute INIT_2A of inst : label is "628B297C012208198005818462CAFFFFE4BE61E334CE6666662666E4B0618532";
    attribute INIT_2B of inst : label is "0313E9F12009D0013B01A0BC1782F050810039BF0E6984668285606282E8104E";
    attribute INIT_2C of inst : label is "501A324CD7013426A6DEE764990E682091011419BBC4F128F04C0253E3140203";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4051400884880A236194C00021242";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "41B8EC4AA2AD486001D143C12AA4D844AACB2AE821D1A40B2038D61526A91036";
    attribute INIT_31 of inst : label is "36B2E45EBAF12E9D120D795EEBC4817B42440503FFB2AA1544889BCB2798AAF6";
    attribute INIT_32 of inst : label is "E0AD2BD569B75F6290DE797AEF3C49EEF3C4BFFBEABCD3617A74D8179A57ABCD";
    attribute INIT_33 of inst : label is "2DB9C2BC063166162C542507A2F1A9950DAA659276218A204408ACFD05EABD36";
    attribute INIT_34 of inst : label is "06082E08905DA82ED4971418EE3D14F153332C1A08A8D21A002A6A294AA8A8C7";
    attribute INIT_35 of inst : label is "45D08D6564FFFFFFFFFA10C48539108C4E2BC86A255D9800429485BA0B830497";
    attribute INIT_36 of inst : label is "82276792C9422AEA5B4014BCE47704D6E4FEDEE257E4874CE1FBB8FE4E031701";
    attribute INIT_37 of inst : label is "D6BC2436496B456CFA64C183264C19026080902601EB9080B800064D2C8B0D38";
    attribute INIT_38 of inst : label is "12D50B321164B46459542C5A4AAAE227B2BCBDAA6A36FA28032C225912E790B1";
    attribute INIT_39 of inst : label is "CE6666662746E6666662746F7F1678665620156D18BBFFE40412D0B446CB2D0B";
    attribute INIT_3A of inst : label is "628B297C012208198005818462CAFFFFE4BE61E334CE6666662666E4B0618532";
    attribute INIT_3B of inst : label is "0313E9F12009D0013B01A0BC1782F050810039BF0E6984668285606282E8104E";
    attribute INIT_3C of inst : label is "501A324CD7013426A6DEE764990E682091011419BBC4F128F04C0253E3140203";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4051400884880A236194C00021242";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "69DEFE7D0761AEB1BDB97FC3FA8EB6CFEA8A3AB1C1D9F375B6AA5B65C7EFC8BF";
    attribute INIT_01 of inst : label is "9B51BCD40ED9B4689B576DC83B66D56F51926DED5EEE0A0000CCDBF5BAF9AAFB";
    attribute INIT_02 of inst : label is "0AEDE9076CD805F6857C6DD03E366C83E366D52D40F8D9B9D1A26D5F1BD20F8D";
    attribute INIT_03 of inst : label is "A75162D318A1FDE53316F5F3D6B8F43FA0FD0D87C5E0A06528852AFD0740FD9B";
    attribute INIT_04 of inst : label is "52977AA12CF4377A1B3D50D8FA3C56F15444054030EED9B3962B6C616553AE45";
    attribute INIT_05 of inst : label is "156F95416CFFFFFFFFF9C74A71D9CE342F87465E7055954A1294A5AD9EA86BBD";
    attribute INIT_06 of inst : label is "F236FBFF6F3264496E6053AFB8F5408424FEDEA1C2AAFF0CE050ACFE24121555";
    attribute INIT_07 of inst : label is "81161E5B6DD58868F80008102040002004091020082240408028EC7B3C9C4DBC";
    attribute INIT_08 of inst : label is "83648D3BB1B5F6761D92346E7AAAF337DB48C610CEFFFBA653F6FBEDBFE0D8F9";
    attribute INIT_09 of inst : label is "77FF9E781E1E7FF9E781E1E19098007878280295E1BFFFEAACBD79F6E4ED7D8D";
    attribute INIT_0A of inst : label is "0A22097E67660A19C2088BF66882FFFF809819990890006187E1E1FF69FE1CEB";
    attribute INIT_0B of inst : label is "5DCAB5550755F0EAAEBEA6A99532A62176EA116A73B85C322102A1310AB76EC2";
    attribute INIT_0C of inst : label is "E59F9EF767655F7B74342586ECEB88AADF9AACD0AFE4F7C348B620A520388220";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE18882008FEEAB62111D75B0A1BE4";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "69DEFE7D0761AEB1BDB97FC3FA8EB6CFEA8A3AB1C1D9F375B6AA5B65C7EFC8BF";
    attribute INIT_11 of inst : label is "9B51BCD40ED9B4689B576DC83B66D56F51926DED5EEE0A0000CCDBF5BAF9AAFB";
    attribute INIT_12 of inst : label is "0AEDE9076CD805F6857C6DD03E366C83E366D52D40F8D9B9D1A26D5F1BD20F8D";
    attribute INIT_13 of inst : label is "A75162D318A1FDE53316F5F3D6B8F43FA0FD0D87C5E0A06528852AFD0740FD9B";
    attribute INIT_14 of inst : label is "52977AA12CF4377A1B3D50D8FA3C56F15444054030EED9B3962B6C616553AE45";
    attribute INIT_15 of inst : label is "156F95416CFFFFFFFFF9C74A71D9CE342F87465E7055954A1294A5AD9EA86BBD";
    attribute INIT_16 of inst : label is "F236FBFF6F3264496E6053AFB8F5408424FEDEA1C2AAFF0CE050ACFE24121555";
    attribute INIT_17 of inst : label is "81161E5B6DD58868F80008102040002004091020082240408028EC7B3C9C4DBC";
    attribute INIT_18 of inst : label is "83648D3BB1B5F6761D92346E7AAAF337DB48C610CEFFFBA653F6FBEDBFE0D8F9";
    attribute INIT_19 of inst : label is "77FF9E781E1E7FF9E781E1E19098007878280295E1BFFFEAACBD79F6E4ED7D8D";
    attribute INIT_1A of inst : label is "0A22097E67660A19C2088BF66882FFFF809819990890006187E1E1FF69FE1CEB";
    attribute INIT_1B of inst : label is "5DCAB5550755F0EAAEBEA6A99532A62176EA116A73B85C322102A1310AB76EC2";
    attribute INIT_1C of inst : label is "E59F9EF767655F7B74342586ECEB88AADF9AACD0AFE4F7C348B620A520388220";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE18882008FEEAB62111D75B0A1BE4";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "69DEFE7D0761AEB1BDB97FC3FA8EB6CFEA8A3AB1C1D9F375B6AA5B65C7EFC8BF";
    attribute INIT_21 of inst : label is "9B51BCD40ED9B4689B576DC83B66D56F51926DED5EEE0A0000CCDBF5BAF9AAFB";
    attribute INIT_22 of inst : label is "0AEDE9076CD805F6857C6DD03E366C83E366D52D40F8D9B9D1A26D5F1BD20F8D";
    attribute INIT_23 of inst : label is "A75162D318A1FDE53316F5F3D6B8F43FA0FD0D87C5E0A06528852AFD0740FD9B";
    attribute INIT_24 of inst : label is "52977AA12CF4377A1B3D50D8FA3C56F15444054030EED9B3962B6C616553AE45";
    attribute INIT_25 of inst : label is "156F95416CFFFFFFFFF9C74A71D9CE342F87465E7055954A1294A5AD9EA86BBD";
    attribute INIT_26 of inst : label is "F236FBFF6F3264496E6053AFB8F5408424FEDEA1C2AAFF0CE050ACFE24121555";
    attribute INIT_27 of inst : label is "81161E5B6DD58868F80008102040002004091020082240408028EC7B3C9C4DBC";
    attribute INIT_28 of inst : label is "83648D3BB1B5F6761D92346E7AAAF337DB48C610CEFFFBA653F6FBEDBFE0D8F9";
    attribute INIT_29 of inst : label is "77FF9E781E1E7FF9E781E1E19098007878280295E1BFFFEAACBD79F6E4ED7D8D";
    attribute INIT_2A of inst : label is "0A22097E67660A19C2088BF66882FFFF809819990890006187E1E1FF69FE1CEB";
    attribute INIT_2B of inst : label is "5DCAB5550755F0EAAEBEA6A99532A62176EA116A73B85C322102A1310AB76EC2";
    attribute INIT_2C of inst : label is "E59F9EF767655F7B74342586ECEB88AADF9AACD0AFE4F7C348B620A520388220";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE18882008FEEAB62111D75B0A1BE4";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "69DEFE7D0761AEB1BDB97FC3FA8EB6CFEA8A3AB1C1D9F375B6AA5B65C7EFC8BF";
    attribute INIT_31 of inst : label is "9B51BCD40ED9B4689B576DC83B66D56F51926DED5EEE0A0000CCDBF5BAF9AAFB";
    attribute INIT_32 of inst : label is "0AEDE9076CD805F6857C6DD03E366C83E366D52D40F8D9B9D1A26D5F1BD20F8D";
    attribute INIT_33 of inst : label is "A75162D318A1FDE53316F5F3D6B8F43FA0FD0D87C5E0A06528852AFD0740FD9B";
    attribute INIT_34 of inst : label is "52977AA12CF4377A1B3D50D8FA3C56F15444054030EED9B3962B6C616553AE45";
    attribute INIT_35 of inst : label is "156F95416CFFFFFFFFF9C74A71D9CE342F87465E7055954A1294A5AD9EA86BBD";
    attribute INIT_36 of inst : label is "F236FBFF6F3264496E6053AFB8F5408424FEDEA1C2AAFF0CE050ACFE24121555";
    attribute INIT_37 of inst : label is "81161E5B6DD58868F80008102040002004091020082240408028EC7B3C9C4DBC";
    attribute INIT_38 of inst : label is "83648D3BB1B5F6761D92346E7AAAF337DB48C610CEFFFBA653F6FBEDBFE0D8F9";
    attribute INIT_39 of inst : label is "77FF9E781E1E7FF9E781E1E19098007878280295E1BFFFEAACBD79F6E4ED7D8D";
    attribute INIT_3A of inst : label is "0A22097E67660A19C2088BF66882FFFF809819990890006187E1E1FF69FE1CEB";
    attribute INIT_3B of inst : label is "5DCAB5550755F0EAAEBEA6A99532A62176EA116A73B85C322102A1310AB76EC2";
    attribute INIT_3C of inst : label is "E59F9EF767655F7B74342586ECEB88AADF9AACD0AFE4F7C348B620A520388220";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE18882008FEEAB62111D75B0A1BE4";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "3A4C7F3F7FDDEEF16AFDE036DE0726A279BD9E7CA59EB93592CC7D298AD2584B";
    attribute INIT_01 of inst : label is "9B14F995AC59B4A94BD62CEAB166C47ED09667885FD5367FEC0A6FF59080E2BB";
    attribute INIT_02 of inst : label is "5AC5CD562CD88F8CA76C2CD3B6166EFB6166D47E4ED859B4D2A52DDB0B9BED85";
    attribute INIT_03 of inst : label is "B35362DA944B88B87ED69DA3E638F01F80FC0587C6252B244488B4FF565AD59B";
    attribute INIT_04 of inst : label is "44156288AAC635631AB15654DA337CC33000651334767B1F9727FF5170C14F4D";
    attribute INIT_05 of inst : label is "066954F52CFFFFFFFFF8F1043D008780CF830C88404C1B5AD6B9CD8D18A30AB1";
    attribute INIT_06 of inst : label is "92894259676BEF6B676CC1893691464B54FEC639232AA28A722D8CFE2412315D";
    attribute INIT_07 of inst : label is "CFA2F3CB2CFFCCF4FE0C183060C103060C183060815D5A9080B0A86EA8BC01A8";
    attribute INIT_08 of inst : label is "BB71DDBBC1B067F6FDF7766E2FE2B28FD9086A9BE86DB3ADC0974DACC9BEDCF8";
    attribute INIT_09 of inst : label is "A82D61FFB4CB02D61FFB4CB2828A007F804A02498386FFFA284F6C6639EC19ED";
    attribute INIT_0A of inst : label is "E8C7BB064F41A69FBAA68A0651EEFFFF8240060452282D0078552A82D607E756";
    attribute INIT_0B of inst : label is "54D23D3C415D382BA725058F91F23E4176EC35E37077B1CEFA4550F202376EB9";
    attribute INIT_0C of inst : label is "F59348E6DC3657F6BB736582C653C9885896FECD8FA4F464490640013994C46B";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC220A00004E9AA8E5B95724998CB25";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "3A4C7F3F7FDDEEF16AFDE036DE0726A279BD9E7CA59EB93592CC7D298AD2584B";
    attribute INIT_11 of inst : label is "9B14F995AC59B4A94BD62CEAB166C47ED09667885FD5367FEC0A6FF59080E2BB";
    attribute INIT_12 of inst : label is "5AC5CD562CD88F8CA76C2CD3B6166EFB6166D47E4ED859B4D2A52DDB0B9BED85";
    attribute INIT_13 of inst : label is "B35362DA944B88B87ED69DA3E638F01F80FC0587C6252B244488B4FF565AD59B";
    attribute INIT_14 of inst : label is "44156288AAC635631AB15654DA337CC33000651334767B1F9727FF5170C14F4D";
    attribute INIT_15 of inst : label is "066954F52CFFFFFFFFF8F1043D008780CF830C88404C1B5AD6B9CD8D18A30AB1";
    attribute INIT_16 of inst : label is "92894259676BEF6B676CC1893691464B54FEC639232AA28A722D8CFE2412315D";
    attribute INIT_17 of inst : label is "CFA2F3CB2CFFCCF4FE0C183060C103060C183060815D5A9080B0A86EA8BC01A8";
    attribute INIT_18 of inst : label is "BB71DDBBC1B067F6FDF7766E2FE2B28FD9086A9BE86DB3ADC0974DACC9BEDCF8";
    attribute INIT_19 of inst : label is "A82D61FFB4CB02D61FFB4CB2828A007F804A02498386FFFA284F6C6639EC19ED";
    attribute INIT_1A of inst : label is "E8C7BB064F41A69FBAA68A0651EEFFFF8240060452282D0078552A82D607E756";
    attribute INIT_1B of inst : label is "54D23D3C415D382BA725058F91F23E4176EC35E37077B1CEFA4550F202376EB9";
    attribute INIT_1C of inst : label is "F59348E6DC3657F6BB736582C653C9885896FECD8FA4F464490640013994C46B";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC220A00004E9AA8E5B95724998CB25";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "3A4C7F3F7FDDEEF16AFDE036DE0726A279BD9E7CA59EB93592CC7D298AD2584B";
    attribute INIT_21 of inst : label is "9B14F995AC59B4A94BD62CEAB166C47ED09667885FD5367FEC0A6FF59080E2BB";
    attribute INIT_22 of inst : label is "5AC5CD562CD88F8CA76C2CD3B6166EFB6166D47E4ED859B4D2A52DDB0B9BED85";
    attribute INIT_23 of inst : label is "B35362DA944B88B87ED69DA3E638F01F80FC0587C6252B244488B4FF565AD59B";
    attribute INIT_24 of inst : label is "44156288AAC635631AB15654DA337CC33000651334767B1F9727FF5170C14F4D";
    attribute INIT_25 of inst : label is "066954F52CFFFFFFFFF8F1043D008780CF830C88404C1B5AD6B9CD8D18A30AB1";
    attribute INIT_26 of inst : label is "92894259676BEF6B676CC1893691464B54FEC639232AA28A722D8CFE2412315D";
    attribute INIT_27 of inst : label is "CFA2F3CB2CFFCCF4FE0C183060C103060C183060815D5A9080B0A86EA8BC01A8";
    attribute INIT_28 of inst : label is "BB71DDBBC1B067F6FDF7766E2FE2B28FD9086A9BE86DB3ADC0974DACC9BEDCF8";
    attribute INIT_29 of inst : label is "A82D61FFB4CB02D61FFB4CB2828A007F804A02498386FFFA284F6C6639EC19ED";
    attribute INIT_2A of inst : label is "E8C7BB064F41A69FBAA68A0651EEFFFF8240060452282D0078552A82D607E756";
    attribute INIT_2B of inst : label is "54D23D3C415D382BA725058F91F23E4176EC35E37077B1CEFA4550F202376EB9";
    attribute INIT_2C of inst : label is "F59348E6DC3657F6BB736582C653C9885896FECD8FA4F464490640013994C46B";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC220A00004E9AA8E5B95724998CB25";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "3A4C7F3F7FDDEEF16AFDE036DE0726A279BD9E7CA59EB93592CC7D298AD2584B";
    attribute INIT_31 of inst : label is "9B14F995AC59B4A94BD62CEAB166C47ED09667885FD5367FEC0A6FF59080E2BB";
    attribute INIT_32 of inst : label is "5AC5CD562CD88F8CA76C2CD3B6166EFB6166D47E4ED859B4D2A52DDB0B9BED85";
    attribute INIT_33 of inst : label is "B35362DA944B88B87ED69DA3E638F01F80FC0587C6252B244488B4FF565AD59B";
    attribute INIT_34 of inst : label is "44156288AAC635631AB15654DA337CC33000651334767B1F9727FF5170C14F4D";
    attribute INIT_35 of inst : label is "066954F52CFFFFFFFFF8F1043D008780CF830C88404C1B5AD6B9CD8D18A30AB1";
    attribute INIT_36 of inst : label is "92894259676BEF6B676CC1893691464B54FEC639232AA28A722D8CFE2412315D";
    attribute INIT_37 of inst : label is "CFA2F3CB2CFFCCF4FE0C183060C103060C183060815D5A9080B0A86EA8BC01A8";
    attribute INIT_38 of inst : label is "BB71DDBBC1B067F6FDF7766E2FE2B28FD9086A9BE86DB3ADC0974DACC9BEDCF8";
    attribute INIT_39 of inst : label is "A82D61FFB4CB02D61FFB4CB2828A007F804A02498386FFFA284F6C6639EC19ED";
    attribute INIT_3A of inst : label is "E8C7BB064F41A69FBAA68A0651EEFFFF8240060452282D0078552A82D607E756";
    attribute INIT_3B of inst : label is "54D23D3C415D382BA725058F91F23E4176EC35E37077B1CEFA4550F202376EB9";
    attribute INIT_3C of inst : label is "F59348E6DC3657F6BB736582C653C9885896FECD8FA4F464490640013994C46B";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC220A00004E9AA8E5B95724998CB25";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "2E4A2C79AE492E3219996009BE866E06FAA93EBFA13AB370964459E7AAF6F189";
    attribute INIT_01 of inst : label is "9B15B175EFD9B58B5BF6CF4FBF66C02C540015CD5000106AB8C95B5090006811";
    attribute INIT_02 of inst : label is "1ED9B9F7ECDA858BAF6D8F57BED66CFBED66D02C5EFB59BF562D6FDB6373EFB5";
    attribute INIT_03 of inst : label is "ACD372DDE069ECAC3CB695B2D634E41F20F9075EC7144188312692FC7D5EFD9B";
    attribute INIT_04 of inst : label is "81196302B0C4B9627C318114AE33B4C338000A0504EC589F000B6D6561873D6D";
    attribute INIT_05 of inst : label is "0671540509FFFFFFFFFA020080201008000C00A00419038CE390C78E18C08C31";
    attribute INIT_06 of inst : label is "BE4508D92F32E4496E6A438AB091910453FEE63A4A2044FD28818BFEC4623959";
    attribute INIT_07 of inst : label is "9127269B6DD18940F80400100040800200080020408800324A52E270C9B8018C";
    attribute INIT_08 of inst : label is "EF60CD1BC7B046B7AD8334EE28E82256894BC832E07D032541B6DAC4D910F8DE";
    attribute INIT_09 of inst : label is "F80000004120FFFFFFFBEDF02D61FF8000001AB58104FFE8A00C3446316C11BD";
    attribute INIT_0A of inst : label is "503024007883023DE4009C404C09FFFFFFFFFFFFFFF800000000007FFFFFFFFF";
    attribute INIT_0B of inst : label is "580E30140150102A02A42488110A2021870917E3CC3615AB094A37A10F3870CA";
    attribute INIT_0C of inst : label is "D4031BD7602956EB604445824CCB5484D85BBC918E91F104914846C26388C120";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF515D500040880AA82A726DB791B17";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "2E4A2C79AE492E3219996009BE866E06FAA93EBFA13AB370964459E7AAF6F189";
    attribute INIT_11 of inst : label is "9B15B175EFD9B58B5BF6CF4FBF66C02C540015CD5000106AB8C95B5090006811";
    attribute INIT_12 of inst : label is "1ED9B9F7ECDA858BAF6D8F57BED66CFBED66D02C5EFB59BF562D6FDB6373EFB5";
    attribute INIT_13 of inst : label is "ACD372DDE069ECAC3CB695B2D634E41F20F9075EC7144188312692FC7D5EFD9B";
    attribute INIT_14 of inst : label is "81196302B0C4B9627C318114AE33B4C338000A0504EC589F000B6D6561873D6D";
    attribute INIT_15 of inst : label is "0671540509FFFFFFFFFA020080201008000C00A00419038CE390C78E18C08C31";
    attribute INIT_16 of inst : label is "BE4508D92F32E4496E6A438AB091910453FEE63A4A2044FD28818BFEC4623959";
    attribute INIT_17 of inst : label is "9127269B6DD18940F80400100040800200080020408800324A52E270C9B8018C";
    attribute INIT_18 of inst : label is "EF60CD1BC7B046B7AD8334EE28E82256894BC832E07D032541B6DAC4D910F8DE";
    attribute INIT_19 of inst : label is "F80000004120FFFFFFFBEDF02D61FF8000001AB58104FFE8A00C3446316C11BD";
    attribute INIT_1A of inst : label is "503024007883023DE4009C404C09FFFFFFFFFFFFFFF800000000007FFFFFFFFF";
    attribute INIT_1B of inst : label is "580E30140150102A02A42488110A2021870917E3CC3615AB094A37A10F3870CA";
    attribute INIT_1C of inst : label is "D4031BD7602956EB604445824CCB5484D85BBC918E91F104914846C26388C120";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF515D500040880AA82A726DB791B17";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "2E4A2C79AE492E3219996009BE866E06FAA93EBFA13AB370964459E7AAF6F189";
    attribute INIT_21 of inst : label is "9B15B175EFD9B58B5BF6CF4FBF66C02C540015CD5000106AB8C95B5090006811";
    attribute INIT_22 of inst : label is "1ED9B9F7ECDA858BAF6D8F57BED66CFBED66D02C5EFB59BF562D6FDB6373EFB5";
    attribute INIT_23 of inst : label is "ACD372DDE069ECAC3CB695B2D634E41F20F9075EC7144188312692FC7D5EFD9B";
    attribute INIT_24 of inst : label is "81196302B0C4B9627C318114AE33B4C338000A0504EC589F000B6D6561873D6D";
    attribute INIT_25 of inst : label is "0671540509FFFFFFFFFA020080201008000C00A00419038CE390C78E18C08C31";
    attribute INIT_26 of inst : label is "BE4508D92F32E4496E6A438AB091910453FEE63A4A2044FD28818BFEC4623959";
    attribute INIT_27 of inst : label is "9127269B6DD18940F80400100040800200080020408800324A52E270C9B8018C";
    attribute INIT_28 of inst : label is "EF60CD1BC7B046B7AD8334EE28E82256894BC832E07D032541B6DAC4D910F8DE";
    attribute INIT_29 of inst : label is "F80000004120FFFFFFFBEDF02D61FF8000001AB58104FFE8A00C3446316C11BD";
    attribute INIT_2A of inst : label is "503024007883023DE4009C404C09FFFFFFFFFFFFFFF800000000007FFFFFFFFF";
    attribute INIT_2B of inst : label is "580E30140150102A02A42488110A2021870917E3CC3615AB094A37A10F3870CA";
    attribute INIT_2C of inst : label is "D4031BD7602956EB604445824CCB5484D85BBC918E91F104914846C26388C120";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF515D500040880AA82A726DB791B17";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "2E4A2C79AE492E3219996009BE866E06FAA93EBFA13AB370964459E7AAF6F189";
    attribute INIT_31 of inst : label is "9B15B175EFD9B58B5BF6CF4FBF66C02C540015CD5000106AB8C95B5090006811";
    attribute INIT_32 of inst : label is "1ED9B9F7ECDA858BAF6D8F57BED66CFBED66D02C5EFB59BF562D6FDB6373EFB5";
    attribute INIT_33 of inst : label is "ACD372DDE069ECAC3CB695B2D634E41F20F9075EC7144188312692FC7D5EFD9B";
    attribute INIT_34 of inst : label is "81196302B0C4B9627C318114AE33B4C338000A0504EC589F000B6D6561873D6D";
    attribute INIT_35 of inst : label is "0671540509FFFFFFFFFA020080201008000C00A00419038CE390C78E18C08C31";
    attribute INIT_36 of inst : label is "BE4508D92F32E4496E6A438AB091910453FEE63A4A2044FD28818BFEC4623959";
    attribute INIT_37 of inst : label is "9127269B6DD18940F80400100040800200080020408800324A52E270C9B8018C";
    attribute INIT_38 of inst : label is "EF60CD1BC7B046B7AD8334EE28E82256894BC832E07D032541B6DAC4D910F8DE";
    attribute INIT_39 of inst : label is "F80000004120FFFFFFFBEDF02D61FF8000001AB58104FFE8A00C3446316C11BD";
    attribute INIT_3A of inst : label is "503024007883023DE4009C404C09FFFFFFFFFFFFFFF800000000007FFFFFFFFF";
    attribute INIT_3B of inst : label is "580E30140150102A02A42488110A2021870917E3CC3615AB094A37A10F3870CA";
    attribute INIT_3C of inst : label is "D4031BD7602956EB604445824CCB5484D85BBC918E91F104914846C26388C120";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF515D500040880AA82A726DB791B17";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "6854D279E65B2F389B996001B8366F76E0AB3839F55AB371B34D596DF2F6E8DB";
    attribute INIT_01 of inst : label is "93142000A81930A14A552C02A064D1083C241572B000296A81ABB711BD0E0143";
    attribute INIT_02 of inst : label is "4AA580540C980910255D2C02A6864C2A6864D5080A9A1930028529574B00A9A1";
    attribute INIT_03 of inst : label is "80C5EFC501258004B41FA7EACE70C20E10708184C022601C2380D1FCC00A8193";
    attribute INIT_04 of inst : label is "C239A784F34DF8A6DC53C0748A3060C220001F08C0ED5E5105DB6CD3E4936E37";
    attribute INIT_05 of inst : label is "1CF626C593FFFFFFFFF808080201004080100800408810429000059E69E11C53";
    attribute INIT_06 of inst : label is "DEEC104B6F3A65596E74439AB393D22C4BFFC66DC6704DBBAC81DBFE442253B1";
    attribute INIT_07 of inst : label is "B56484934D59B353F8040800004080020400002040291281B11D316102D061C3";
    attribute INIT_08 of inst : label is "0B482DDB85B094B42D20B76F4A816AEE1290DA7661B66AE2012492C952749A9A";
    attribute INIT_09 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFB0B5254005FFE877967494516C252D";
    attribute INIT_0A of inst : label is "F8862001FC16064AE802AC218188FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000";
    attribute INIT_0B of inst : label is "B022700006B000D600583A9A334E69939B1245A74915B30B548180AC9F79B15E";
    attribute INIT_0C of inst : label is "9E6B999600E1864028547586CCDB0880D83199219C0BF0000000070805000203";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2A2A000A8A9C19424526DB485B0C";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "6854D279E65B2F389B996001B8366F76E0AB3839F55AB371B34D596DF2F6E8DB";
    attribute INIT_11 of inst : label is "93142000A81930A14A552C02A064D1083C241572B000296A81ABB711BD0E0143";
    attribute INIT_12 of inst : label is "4AA580540C980910255D2C02A6864C2A6864D5080A9A1930028529574B00A9A1";
    attribute INIT_13 of inst : label is "80C5EFC501258004B41FA7EACE70C20E10708184C022601C2380D1FCC00A8193";
    attribute INIT_14 of inst : label is "C239A784F34DF8A6DC53C0748A3060C220001F08C0ED5E5105DB6CD3E4936E37";
    attribute INIT_15 of inst : label is "1CF626C593FFFFFFFFF808080201004080100800408810429000059E69E11C53";
    attribute INIT_16 of inst : label is "DEEC104B6F3A65596E74439AB393D22C4BFFC66DC6704DBBAC81DBFE442253B1";
    attribute INIT_17 of inst : label is "B56484934D59B353F8040800004080020400002040291281B11D316102D061C3";
    attribute INIT_18 of inst : label is "0B482DDB85B094B42D20B76F4A816AEE1290DA7661B66AE2012492C952749A9A";
    attribute INIT_19 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFB0B5254005FFE877967494516C252D";
    attribute INIT_1A of inst : label is "F8862001FC16064AE802AC218188FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000";
    attribute INIT_1B of inst : label is "B022700006B000D600583A9A334E69939B1245A74915B30B548180AC9F79B15E";
    attribute INIT_1C of inst : label is "9E6B999600E1864028547586CCDB0880D83199219C0BF0000000070805000203";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2A2A000A8A9C19424526DB485B0C";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "6854D279E65B2F389B996001B8366F76E0AB3839F55AB371B34D596DF2F6E8DB";
    attribute INIT_21 of inst : label is "93142000A81930A14A552C02A064D1083C241572B000296A81ABB711BD0E0143";
    attribute INIT_22 of inst : label is "4AA580540C980910255D2C02A6864C2A6864D5080A9A1930028529574B00A9A1";
    attribute INIT_23 of inst : label is "80C5EFC501258004B41FA7EACE70C20E10708184C022601C2380D1FCC00A8193";
    attribute INIT_24 of inst : label is "C239A784F34DF8A6DC53C0748A3060C220001F08C0ED5E5105DB6CD3E4936E37";
    attribute INIT_25 of inst : label is "1CF626C593FFFFFFFFF808080201004080100800408810429000059E69E11C53";
    attribute INIT_26 of inst : label is "DEEC104B6F3A65596E74439AB393D22C4BFFC66DC6704DBBAC81DBFE442253B1";
    attribute INIT_27 of inst : label is "B56484934D59B353F8040800004080020400002040291281B11D316102D061C3";
    attribute INIT_28 of inst : label is "0B482DDB85B094B42D20B76F4A816AEE1290DA7661B66AE2012492C952749A9A";
    attribute INIT_29 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFB0B5254005FFE877967494516C252D";
    attribute INIT_2A of inst : label is "F8862001FC16064AE802AC218188FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000";
    attribute INIT_2B of inst : label is "B022700006B000D600583A9A334E69939B1245A74915B30B548180AC9F79B15E";
    attribute INIT_2C of inst : label is "9E6B999600E1864028547586CCDB0880D83199219C0BF0000000070805000203";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2A2A000A8A9C19424526DB485B0C";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "6854D279E65B2F389B996001B8366F76E0AB3839F55AB371B34D596DF2F6E8DB";
    attribute INIT_31 of inst : label is "93142000A81930A14A552C02A064D1083C241572B000296A81ABB711BD0E0143";
    attribute INIT_32 of inst : label is "4AA580540C980910255D2C02A6864C2A6864D5080A9A1930028529574B00A9A1";
    attribute INIT_33 of inst : label is "80C5EFC501258004B41FA7EACE70C20E10708184C022601C2380D1FCC00A8193";
    attribute INIT_34 of inst : label is "C239A784F34DF8A6DC53C0748A3060C220001F08C0ED5E5105DB6CD3E4936E37";
    attribute INIT_35 of inst : label is "1CF626C593FFFFFFFFF808080201004080100800408810429000059E69E11C53";
    attribute INIT_36 of inst : label is "DEEC104B6F3A65596E74439AB393D22C4BFFC66DC6704DBBAC81DBFE442253B1";
    attribute INIT_37 of inst : label is "B56484934D59B353F8040800004080020400002040291281B11D316102D061C3";
    attribute INIT_38 of inst : label is "0B482DDB85B094B42D20B76F4A816AEE1290DA7661B66AE2012492C952749A9A";
    attribute INIT_39 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFB0B5254005FFE877967494516C252D";
    attribute INIT_3A of inst : label is "F8862001FC16064AE802AC218188FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000";
    attribute INIT_3B of inst : label is "B022700006B000D600583A9A334E69939B1245A74915B30B548180AC9F79B15E";
    attribute INIT_3C of inst : label is "9E6B999600E1864028547586CCDB0880D83199219C0BF0000000070805000203";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2A2A000A8A9C19424526DB485B0C";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "789E7F6B80C16DB9C85D60059A076DA6E80EBA30895CBB65BDEC5B218AC6F89B";
    attribute INIT_01 of inst : label is "CB44B2034EDCB3660BA76C253B72D42CCDB645FD500026D567098325BAC5A24B";
    attribute INIT_02 of inst : label is "34ED84A76E5A0D901A786C0D3C372E53C372C42C34F0DCB80D982E9E1B094F0D";
    attribute INIT_03 of inst : label is "96C366C21129A00532579DE2E6141800C00602A905A823044088A4FF6034EDCB";
    attribute INIT_04 of inst : label is "444560880AC34561A2B04414383300C000006113106459119203EF4D76D90E2D";
    attribute INIT_05 of inst : label is "1C0F18730EFFFFFFFFFBF790FDF21FB90FEF90FC8777239C61084CC118222230";
    attribute INIT_06 of inst : label is "E77298DB6D720C4B6D7541813E90460714FF4B17A2137D99F27C86FE884650E4";
    attribute INIT_07 of inst : label is "C69716DB6DEDCC24FD8E1E3878A162C70F1C3C50B08DB2E5077FDA7741846181";
    attribute INIT_08 of inst : label is "8165840B08B256160596102C25A262665B2C6388E9FD4B2C40B6D96DD9565858";
    attribute INIT_09 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFE4327DE181FFF3DACB5E57302C9585";
    attribute INIT_0A of inst : label is "A8C39107376E0000F908F67310E4FFFF80000000000000000000000000000000";
    attribute INIT_0B of inst : label is "EC12040407E402FC813E6F8190320740448EC1A139840D233604A43A0E0448F3";
    attribute INIT_0C of inst : label is "3B4BDB36FCED4617871F0586C6437A825CDE601C8134F7CDF37CC0F7FAF904A0";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B27321A388322DBC80B36";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "789E7F6B80C16DB9C85D60059A076DA6E80EBA30895CBB65BDEC5B218AC6F89B";
    attribute INIT_11 of inst : label is "CB44B2034EDCB3660BA76C253B72D42CCDB645FD500026D567098325BAC5A24B";
    attribute INIT_12 of inst : label is "34ED84A76E5A0D901A786C0D3C372E53C372C42C34F0DCB80D982E9E1B094F0D";
    attribute INIT_13 of inst : label is "96C366C21129A00532579DE2E6141800C00602A905A823044088A4FF6034EDCB";
    attribute INIT_14 of inst : label is "444560880AC34561A2B04414383300C000006113106459119203EF4D76D90E2D";
    attribute INIT_15 of inst : label is "1C0F18730EFFFFFFFFFBF790FDF21FB90FEF90FC8777239C61084CC118222230";
    attribute INIT_16 of inst : label is "E77298DB6D720C4B6D7541813E90460714FF4B17A2137D99F27C86FE884650E4";
    attribute INIT_17 of inst : label is "C69716DB6DEDCC24FD8E1E3878A162C70F1C3C50B08DB2E5077FDA7741846181";
    attribute INIT_18 of inst : label is "8165840B08B256160596102C25A262665B2C6388E9FD4B2C40B6D96DD9565858";
    attribute INIT_19 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFE4327DE181FFF3DACB5E57302C9585";
    attribute INIT_1A of inst : label is "A8C39107376E0000F908F67310E4FFFF80000000000000000000000000000000";
    attribute INIT_1B of inst : label is "EC12040407E402FC813E6F8190320740448EC1A139840D233604A43A0E0448F3";
    attribute INIT_1C of inst : label is "3B4BDB36FCED4617871F0586C6437A825CDE601C8134F7CDF37CC0F7FAF904A0";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B27321A388322DBC80B36";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "789E7F6B80C16DB9C85D60059A076DA6E80EBA30895CBB65BDEC5B218AC6F89B";
    attribute INIT_21 of inst : label is "CB44B2034EDCB3660BA76C253B72D42CCDB645FD500026D567098325BAC5A24B";
    attribute INIT_22 of inst : label is "34ED84A76E5A0D901A786C0D3C372E53C372C42C34F0DCB80D982E9E1B094F0D";
    attribute INIT_23 of inst : label is "96C366C21129A00532579DE2E6141800C00602A905A823044088A4FF6034EDCB";
    attribute INIT_24 of inst : label is "444560880AC34561A2B04414383300C000006113106459119203EF4D76D90E2D";
    attribute INIT_25 of inst : label is "1C0F18730EFFFFFFFFFBF790FDF21FB90FEF90FC8777239C61084CC118222230";
    attribute INIT_26 of inst : label is "E77298DB6D720C4B6D7541813E90460714FF4B17A2137D99F27C86FE884650E4";
    attribute INIT_27 of inst : label is "C69716DB6DEDCC24FD8E1E3878A162C70F1C3C50B08DB2E5077FDA7741846181";
    attribute INIT_28 of inst : label is "8165840B08B256160596102C25A262665B2C6388E9FD4B2C40B6D96DD9565858";
    attribute INIT_29 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFE4327DE181FFF3DACB5E57302C9585";
    attribute INIT_2A of inst : label is "A8C39107376E0000F908F67310E4FFFF80000000000000000000000000000000";
    attribute INIT_2B of inst : label is "EC12040407E402FC813E6F8190320740448EC1A139840D233604A43A0E0448F3";
    attribute INIT_2C of inst : label is "3B4BDB36FCED4617871F0586C6437A825CDE601C8134F7CDF37CC0F7FAF904A0";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B27321A388322DBC80B36";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "789E7F6B80C16DB9C85D60059A076DA6E80EBA30895CBB65BDEC5B218AC6F89B";
    attribute INIT_31 of inst : label is "CB44B2034EDCB3660BA76C253B72D42CCDB645FD500026D567098325BAC5A24B";
    attribute INIT_32 of inst : label is "34ED84A76E5A0D901A786C0D3C372E53C372C42C34F0DCB80D982E9E1B094F0D";
    attribute INIT_33 of inst : label is "96C366C21129A00532579DE2E6141800C00602A905A823044088A4FF6034EDCB";
    attribute INIT_34 of inst : label is "444560880AC34561A2B04414383300C000006113106459119203EF4D76D90E2D";
    attribute INIT_35 of inst : label is "1C0F18730EFFFFFFFFFBF790FDF21FB90FEF90FC8777239C61084CC118222230";
    attribute INIT_36 of inst : label is "E77298DB6D720C4B6D7541813E90460714FF4B17A2137D99F27C86FE884650E4";
    attribute INIT_37 of inst : label is "C69716DB6DEDCC24FD8E1E3878A162C70F1C3C50B08DB2E5077FDA7741846181";
    attribute INIT_38 of inst : label is "8165840B08B256160596102C25A262665B2C6388E9FD4B2C40B6D96DD9565858";
    attribute INIT_39 of inst : label is "0000000000007FFFFFFBEDF7FFFFFFFFFFE4327DE181FFF3DACB5E57302C9585";
    attribute INIT_3A of inst : label is "A8C39107376E0000F908F67310E4FFFF80000000000000000000000000000000";
    attribute INIT_3B of inst : label is "EC12040407E402FC813E6F8190320740448EC1A139840D233604A43A0E0448F3";
    attribute INIT_3C of inst : label is "3B4BDB36FCED4617871F0586C6437A825CDE601C8134F7CDF37CC0F7FAF904A0";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B27321A388322DBC80B36";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "3914132BA2C8659FC9CD2004B0632582400A9018894C992C9D8849248A426889";
    attribute INIT_01 of inst : label is "D9AE920BE48D9BB719F2443792367FE4CFDFC4FC00002D956719936C98410459";
    attribute INIT_02 of inst : label is "BE4886F246CF5C907F28442F9423677942367BE4BE508D982EDC67CA110DE508";
    attribute INIT_03 of inst : label is "964126473B38914717D3DCE246181008A04402A981C4606C0D8120FEA0BE48D9";
    attribute INIT_04 of inst : label is "C28E61851CC00E600730C298183054C15400570810644B10DE89E44F3E792624";
    attribute INIT_05 of inst : label is "1C1F94204AFFFFFFFFF8000800010000800008004000125296B5ACC3D86147B0";
    attribute INIT_06 of inst : label is "E264984925722C43273541879A90C2C220FE4215C21B7909806882FE040050EC";
    attribute INIT_07 of inst : label is "8A02734924EC8820FA81000008100140A000840A015FB0E587AFDC3340847C80";
    attribute INIT_08 of inst : label is "83218C190192D2320C86306467044666C9244700E9EF490E40924D648B4AC8C8";
    attribute INIT_09 of inst : label is "FFFFFFFFFFFF80000004120800000000006432D8E119FFF7D8DB5AD36064B48C";
    attribute INIT_0A of inst : label is "B88100383C0E0020D908F2700040FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0B of inst : label is "E4820C0407EC02FD803E2FC718EB1C00E5CEC12111840523F400A0200E0E5C90";
    attribute INIT_0C of inst : label is "2B89CB33BCF6421D823A04824649BA8ECC1A20088100F00401004000000086A0";
    attribute INIT_0D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B67321411010249C81906";
    attribute INIT_0E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_10 of inst : label is "3914132BA2C8659FC9CD2004B0632582400A9018894C992C9D8849248A426889";
    attribute INIT_11 of inst : label is "D9AE920BE48D9BB719F2443792367FE4CFDFC4FC00002D956719936C98410459";
    attribute INIT_12 of inst : label is "BE4886F246CF5C907F28442F9423677942367BE4BE508D982EDC67CA110DE508";
    attribute INIT_13 of inst : label is "964126473B38914717D3DCE246181008A04402A981C4606C0D8120FEA0BE48D9";
    attribute INIT_14 of inst : label is "C28E61851CC00E600730C298183054C15400570810644B10DE89E44F3E792624";
    attribute INIT_15 of inst : label is "1C1F94204AFFFFFFFFF8000800010000800008004000125296B5ACC3D86147B0";
    attribute INIT_16 of inst : label is "E264984925722C43273541879A90C2C220FE4215C21B7909806882FE040050EC";
    attribute INIT_17 of inst : label is "8A02734924EC8820FA81000008100140A000840A015FB0E587AFDC3340847C80";
    attribute INIT_18 of inst : label is "83218C190192D2320C86306467044666C9244700E9EF490E40924D648B4AC8C8";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFF80000004120800000000006432D8E119FFF7D8DB5AD36064B48C";
    attribute INIT_1A of inst : label is "B88100383C0E0020D908F2700040FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1B of inst : label is "E4820C0407EC02FD803E2FC718EB1C00E5CEC12111840523F400A0200E0E5C90";
    attribute INIT_1C of inst : label is "2B89CB33BCF6421D823A04824649BA8ECC1A20088100F00401004000000086A0";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B67321411010249C81906";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "3914132BA2C8659FC9CD2004B0632582400A9018894C992C9D8849248A426889";
    attribute INIT_21 of inst : label is "D9AE920BE48D9BB719F2443792367FE4CFDFC4FC00002D956719936C98410459";
    attribute INIT_22 of inst : label is "BE4886F246CF5C907F28442F9423677942367BE4BE508D982EDC67CA110DE508";
    attribute INIT_23 of inst : label is "964126473B38914717D3DCE246181008A04402A981C4606C0D8120FEA0BE48D9";
    attribute INIT_24 of inst : label is "C28E61851CC00E600730C298183054C15400570810644B10DE89E44F3E792624";
    attribute INIT_25 of inst : label is "1C1F94204AFFFFFFFFF8000800010000800008004000125296B5ACC3D86147B0";
    attribute INIT_26 of inst : label is "E264984925722C43273541879A90C2C220FE4215C21B7909806882FE040050EC";
    attribute INIT_27 of inst : label is "8A02734924EC8820FA81000008100140A000840A015FB0E587AFDC3340847C80";
    attribute INIT_28 of inst : label is "83218C190192D2320C86306467044666C9244700E9EF490E40924D648B4AC8C8";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFF80000004120800000000006432D8E119FFF7D8DB5AD36064B48C";
    attribute INIT_2A of inst : label is "B88100383C0E0020D908F2700040FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "E4820C0407EC02FD803E2FC718EB1C00E5CEC12111840523F400A0200E0E5C90";
    attribute INIT_2C of inst : label is "2B89CB33BCF6421D823A04824649BA8ECC1A20088100F00401004000000086A0";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B67321411010249C81906";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "3914132BA2C8659FC9CD2004B0632582400A9018894C992C9D8849248A426889";
    attribute INIT_31 of inst : label is "D9AE920BE48D9BB719F2443792367FE4CFDFC4FC00002D956719936C98410459";
    attribute INIT_32 of inst : label is "BE4886F246CF5C907F28442F9423677942367BE4BE508D982EDC67CA110DE508";
    attribute INIT_33 of inst : label is "964126473B38914717D3DCE246181008A04402A981C4606C0D8120FEA0BE48D9";
    attribute INIT_34 of inst : label is "C28E61851CC00E600730C298183054C15400570810644B10DE89E44F3E792624";
    attribute INIT_35 of inst : label is "1C1F94204AFFFFFFFFF8000800010000800008004000125296B5ACC3D86147B0";
    attribute INIT_36 of inst : label is "E264984925722C43273541879A90C2C220FE4215C21B7909806882FE040050EC";
    attribute INIT_37 of inst : label is "8A02734924EC8820FA81000008100140A000840A015FB0E587AFDC3340847C80";
    attribute INIT_38 of inst : label is "83218C190192D2320C86306467044666C9244700E9EF490E40924D648B4AC8C8";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFF80000004120800000000006432D8E119FFF7D8DB5AD36064B48C";
    attribute INIT_3A of inst : label is "B88100383C0E0020D908F2700040FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "E4820C0407EC02FD803E2FC718EB1C00E5CEC12111840523F400A0200E0E5C90";
    attribute INIT_3C of inst : label is "2B89CB33BCF6421D823A04824649BA8ECC1A20088100F00401004000000086A0";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA2AAA000B67321411010249C81906";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
