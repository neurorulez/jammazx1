-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "499AFFE2175962241C7471D1229333588200FFC000000000010045DFDE5B1307";
    attribute INIT_01 of inst : label is "E200A47A632D4822A05FD7D5FD7954C1015011200A080C5082984B42F08C9B36";
    attribute INIT_02 of inst : label is "1CBC62F1B828904234822D244044A28101128A04027071C38480090A2AB01C7F";
    attribute INIT_03 of inst : label is "E1E96000F40418281240004B4585242CA28E0E181E23CA04108D208348484A55";
    attribute INIT_04 of inst : label is "CDFF700128462F0F44A2452808C5E1C04050988CF1B88A200002383A28800008";
    attribute INIT_05 of inst : label is "5391C33045E18A00707862801C3D029C9016FE13FDE872DFC27FBD53F24DFF75";
    attribute INIT_06 of inst : label is "C0C803404697FF9465105552692C5924912A721CDA2B48D610DC395A4B1BFF37";
    attribute INIT_07 of inst : label is "5FCDD4F158774CC001FC4001790AAC1144DE2A1BC2C5402D561021DA2B48D630";
    attribute INIT_08 of inst : label is "776ABD5FCDC8737776ABD5FCDD4EB2A101409790877FF7BBD5FCD88737FF7BBD";
    attribute INIT_09 of inst : label is "A770608C53FC323E23978CFA9E573737C6357104629FC3F03986D3E1E3822477";
    attribute INIT_0A of inst : label is "224C4437EDFFDDEF74215604108840405E03C07E4C92C00B340309C210012844";
    attribute INIT_0B of inst : label is "CEF670A74C3A8FF905FFD7865436408FFADD13CD5497A5D6AA81706F2A28A901";
    attribute INIT_0C of inst : label is "B005F4D2BBFDAA4C747EC741BF0FD63A858B3FF18EC01F600FC000009DF7171C";
    attribute INIT_0D of inst : label is "C495EFE66B21699FFA6766933FF4CE69B665AD902B96D9A327D273D6CEB6EBCD";
    attribute INIT_0E of inst : label is "A7CE6227FFB8277CF3EEEE64D6B957BDDD9F82CFC422BF5A63EA90892808A3A8";
    attribute INIT_0F of inst : label is "4E4400000001C8820045104000BE78011451001C71E064393F544539F73117FF";
    attribute INIT_10 of inst : label is "482C922F0D525620A64DBDF45D10000000E74514624CA2884957D589268B6E74";
    attribute INIT_11 of inst : label is "2400071A000C42B8008A288019451002AFAA004D16C0089C88000000045F45D1";
    attribute INIT_12 of inst : label is "4AB34074E04559A885A9D428AB86CCFAACC3771342509481081215C680AE3011";
    attribute INIT_13 of inst : label is "4000000000FC3C667FBFAA43121E5CA39320E5C0081002214020A0D360085D1D";
    attribute INIT_14 of inst : label is "D248000325A4C000100804000100924000325B6C001A71EA7FEDFDD49DF8703D";
    attribute INIT_15 of inst : label is "0C000000001B0C000000001B0C00000000021300000DB6180000000000000026";
    attribute INIT_16 of inst : label is "AA0106FBFEAD144005501FB1A4D78A1E6C20E4838A1A6840000000000000001B";
    attribute INIT_17 of inst : label is "C158A528569094AB69CA4826DCB75D222228822228822228822228828280A802";
    attribute INIT_18 of inst : label is "CBDA52A5FB542806FAF13868FE519C6718CE9ABF63E9FB1AFDA180467E90B238";
    attribute INIT_19 of inst : label is "A36DD4A5CCA53AD237BD697840D48DAD6ADAB44081088AFD36ED13095E16ACED";
    attribute INIT_1A of inst : label is "5E6B388E3DAFF10A040837650CEF1506EFF8DEBB295E5295E90B4A54C080FB3D";
    attribute INIT_1B of inst : label is "489C8BFADFABDBD737FD797AF2FF956FAD750204080C33E908BF130D6E58A7B1";
    attribute INIT_1C of inst : label is "206534B1CB5D32D32AD6559CE518CA95A5EB6BD61395A10A46B540810193FB22";
    attribute INIT_1D of inst : label is "4256BC2108468010004081017B052F7D30D6B18C6318D6A18C6B5AD6B5C00810";
    attribute INIT_1E of inst : label is "16BDAEF8FDF6218C6EDAD6A0810204029FC48D1A53A6A533D5ED9BD21095A97B";
    attribute INIT_1F of inst : label is "8AF7B4FF684AB59C293ACE7EFDAD0E579542810804080D37C8341685CCD74EDD";
    attribute INIT_20 of inst : label is "20009CDEC954A996A5AC631DE6BFFF773CC635A9600204081B7BDB9CB348A2C4";
    attribute INIT_21 of inst : label is "82040012C924CA45F30D7EDFB4BF6FDBF6FDBF6FDBF6FDBB4ED3B4ED3F680800";
    attribute INIT_22 of inst : label is "BCE7B94B9BE6F52BCAF640840A040FACA44CB5ACE358C6B18D1F3AAE6DCFDB7A";
    attribute INIT_23 of inst : label is "1EB46640158B58D6A83118E3114909425094248102040126D21619A2672A5EF4";
    attribute INIT_24 of inst : label is "7686812244004000FC93534BDA090C421886314A15B5652E804280020406DDED";
    attribute INIT_25 of inst : label is "D947FCEEFFEBD71FEC31EE20028402000016E88956716995A5285E96AD6B49DE";
    attribute INIT_26 of inst : label is "733FC01D0806F6FE064522BA5D8E5ECE792856D7ACAF4BD21FDF2729CA7C877D";
    attribute INIT_27 of inst : label is "005468005235F0001526000000000000000592D3C09B322501D7DF000000006A";
    attribute INIT_28 of inst : label is "00000000000000000000000000000000000000000000170BCFFFFDF980000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "408808053D9006649566DC88B3841193A64981000000000001000C7E7E320301";
    attribute INIT_01 of inst : label is "CD22F8D3E841ADDB393B3057B301732C933B32B5A5649CB43CFA1027FC1C0BD3";
    attribute INIT_02 of inst : label is "2F10AC5215BD0B3936596C934B2A464D8CF939372456295932496CBBC99679F6";
    attribute INIT_03 of inst : label is "AC8DED84E25DB1396925B4AF49B6B6907197852B08410F62CA4D96732F6F2323";
    attribute INIT_04 of inst : label is "51BF22B29DE409654871671D9C912C9A9B3BDB105214F2E96B2E2B13CBA5ACB8";
    attribute INIT_05 of inst : label is "4866FCD798ADCE99562B73A6559525910100912DFA4B001225BF49284685BF23";
    attribute INIT_06 of inst : label is "0A991565CCED5F38CD24CDDBCE90B6DB59B3B6C013C52765A3915FB3842CBEDA";
    attribute INIT_07 of inst : label is "FFF6921BC185507326206318606CB9599A4CC9320B966D13664CBE13C52764A5";
    attribute INIT_08 of inst : label is "891133FFF6BB004891133FFF692046CE0DDC0606C84891133FFF6BB004891133";
    attribute INIT_09 of inst : label is "B96C5602550504FCCE2259440980BC7F2C2DF37012A81166E046F608C6CDB884";
    attribute INIT_0A of inst : label is "BDB08DB8ADA06DA68694CF733D3FD4D4912724E1ACA00BC0B736E20400000EE3";
    attribute INIT_0B of inst : label is "1280F9A40D40ED03DE9E47BEEEB90997A2CF66147DCC6FC8935E55FE924F3525";
    attribute INIT_0C of inst : label is "E14A895CC854AB9E24A121159047449820C00163356452B229646464533F81BF";
    attribute INIT_0D of inst : label is "D327918C82AB2414A494592829492892C9768A5DB04802CB3A24243A1A262856";
    attribute INIT_0E of inst : label is "AA07EF7030210F19619C2352F2E03E731415AE0AD2F1FFCB6E3EF79C9D996FEF";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000000000F105603EEC1103F7B830";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "C5A00B2C000044B4000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "7F276C6F0B5F93BAD76E1AEC86B52DC38AD3C82C6372CE449C8933CE4BBEF256";
    attribute INIT_13 of inst : label is "600000000003FC1E15552B2674C89112A444881B4B316525C5BCB767ECE93333";
    attribute INIT_14 of inst : label is "F6DA7F27B7FFE4F2592DB64F2592DB77F27B7FFFF60002054DFABD7A39046591";
    attribute INIT_15 of inst : label is "93FFE7F3FFE493FFE7F3FFE493FFE7F209268178FB9FFFFC9249FCB66D27F26F";
    attribute INIT_16 of inst : label is "FBFEAD1440055015501510AF14B91BB07A80BE46A05AC541FFFCFE7FE7F3FFE4";
    attribute INIT_17 of inst : label is "90584402948780086000056D4E16B5228280A28280A28280A28280A802AA0106";
    attribute INIT_18 of inst : label is "C728088C3104280216019C60442539CA5380E229044108E411C040C020835158";
    attribute INIT_19 of inst : label is "33BC286A0C75CE479EFECDCC74DEFE338E6C91028109604041500315258A5925";
    attribute INIT_1A of inst : label is "79D2173DE15AE00004025A2010D42BE643FEEF3B2A4ED7B4417842090000B522";
    attribute INIT_1B of inst : label is "0B2004CA23084319C4611063388C890C67900000000EFA6890DBA91952358EA4";
    attribute INIT_1C of inst : label is "2012A0A92F4015091C6052232A0298C7110A230CC4210E763400000001F7C111";
    attribute INIT_1D of inst : label is "6BA4CE3FEC078840A000000041179436905358C4B5AE6322D6BD8C4B50902000";
    attribute INIT_1E of inst : label is "8698C628CA6B48C7B00D62B800000001C9044BA680BCC4715738D3F8DAEF307F";
    attribute INIT_1F of inst : label is "A4C61028521CC20542619014800878621816045A10000612222C200D82F286C0";
    attribute INIT_20 of inst : label is "00402B514CAA6481E6629405280A408CE219CE76A0080008079E0012F41B1010";
    attribute INIT_21 of inst : label is "C2002017F0AE2C88C911252A55D4A52929421084216B5AD6B5AD6B5AD2940010";
    attribute INIT_22 of inst : label is "11CFE0931FFE3271900002010806FA0ED0A494D631CF7358D789C85312951EB5";
    attribute INIT_23 of inst : label is "0A5077A454E4422920000400004201080010802040000564016A2081222F8020";
    attribute INIT_24 of inst : label is "A9240028002000806289ABE54811000008400010A3284C500000010800071324";
    attribute INIT_25 of inst : label is "84B50928CC618C4420F58C294085020408146C832AB264809E63390E531A8731";
    attribute INIT_26 of inst : label is "1B506BF80202FC8249A287ED75A118D1FC2118A408820108A12977D633A96252";
    attribute INIT_27 of inst : label is "0491F90128FD40000281000000000000000AA06481C289430228A20000000022";
    attribute INIT_28 of inst : label is "000000000000000000000000000000000000000000000F078FFFFDFA00000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "40893101177FF3B62EDC3264CCA05522B100FEC0000000000000052E2E3F0900";
    attribute INIT_01 of inst : label is "3199376E6ADB792CC984A9584A859CB249DCD8E739920834451AB6DBFE0C09F1";
    attribute INIT_02 of inst : label is "5EED6BA5E9EFB68C2DB4EA4D769F2F075A2C9C1D38B5DAD6CD36926C6C77C649";
    attribute INIT_03 of inst : label is "6B66526E93B34ECE8E934F33754DEDE99EAF7B5AF6BEDBEDA70B6D1299D9D3DD";
    attribute INIT_04 of inst : label is "7740D8ECEE6B975A71B1986E6D72EB72F6DC942FA5ED19ACCED25AEC66B33B49";
    attribute INIT_05 of inst : label is "6499E334677A4F91F5DE93E47D69D1AD891A8D3603CCD351A6C0798CB7A340D8";
    attribute INIT_06 of inst : label is "CEF196326FF77DACEDD198DEFF3DDF6D4DE3FB34546399B7B3597EFFCF76FBEE";
    attribute INIT_07 of inst : label is "001B993FE1E5687387A5F39A9A3868F74D330CD0768DD9958070ED546399B7B5";
    attribute INIT_08 of inst : label is "650CCC001B8CD14650CCC001B99226EE6D9C29A3954650CCC001BACD14650CCC";
    attribute INIT_09 of inst : label is "1C16DE50E4FF092BB9A2753406A4DBFF3B6FF3D28727F19CD25B35F832CDB854";
    attribute INIT_0A of inst : label is "64C77748F78C5EA639E70B7669B58484BD20A411C2AD8AF68D96A4C200001C77";
    attribute INIT_0B of inst : label is "1408FE1BA06534FB8E3F98A280A960CA02C344147DE37FE6C45EF77FCB9145CF";
    attribute INIT_0C of inst : label is "E4776DD7AC74F69B370048168F4094B0A1601E19E5467AA33D464646FAFF592B";
    attribute INIT_0D of inst : label is "DD2C566AE4CF012356F50DB246ADEABF6DBE936FEA9E5769ADB7D6EB1A4A093B";
    attribute INIT_0E of inst : label is "AC2F488F8E9908C51C50A59B339C99CA1755B32AD934FE8CB1D5296F6E6C5BD9";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000086465F2AFCF417A4478E";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "48A00A5400026908000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "9567DB470EF2B3E13838A3B858A9B55CB35A20C99983B7866F0C88E78667BC18";
    attribute INIT_13 of inst : label is "60000000000003FE0CE646929F34D7CD31F34D66CED9993B6664E927F32E8E8E";
    attribute INIT_14 of inst : label is "0000360000121B00048121B00048001360000001B61603016FFDFFAB3DC095DD";
    attribute INIT_15 of inst : label is "01B6C301B6C001B6C301B6C001B6C300000000371F0000C16CB0002424036000";
    attribute INIT_16 of inst : label is "14400550155015155550502AFE050FAE9111BAF8000EAEE1B6D86C36C301B6C0";
    attribute INIT_17 of inst : label is "4DBA8C310C608100231CCEC40EEC143802AA0802AA0802AA0802AA0106FBFEAD";
    attribute INIT_18 of inst : label is "095A76420086080A53CA39CA244308421188E618C8430842080840A03C82C4E8";
    attribute INIT_19 of inst : label is "818DA5F8682D292E7184210A465394A72952A90081014AB854DD5A0B4AF5A950";
    attribute INIT_1A of inst : label is "9CE3BA5EBFBDCC0C040750C0027F03FF2EF69CE7ED63988601AFDBC00000B41C";
    attribute INIT_1B of inst : label is "56314FE6D885B000000800210843B88180F40000000AC1AB34C5200F6EDA5430";
    attribute INIT_1C of inst : label is "25235C924E3CD3403C64D312E471000000022108623080162108000000143975";
    attribute INIT_1D of inst : label is "7BE6DFB1CC9722440812000229034E06003084310C40006010084310CC80200C";
    attribute INIT_1E of inst : label is "4796A520286202852FCB7B280000000122E495A3D6101032B6B530F03CC7383F";
    attribute INIT_1F of inst : label is "8C4330B62304012540310CDAF9841CE31942000000001A85809C6EAC3007C308";
    attribute INIT_20 of inst : label is "0000490E486CA016A5AD6FDADF319EEB7EF6F196300800080BB5C124E69AE06B";
    attribute INIT_21 of inst : label is "88100802D72A0DA2201B6F78C5718C6318CE739CE77BDEF5AD6B5AD6B7B02010";
    attribute INIT_22 of inst : label is "00010002139DEC710C6240244802952A45001CA5AD084250850D6E018636D79C";
    attribute INIT_23 of inst : label is "56952F7FEFA2D694AA2118C211096A5294B5AC000000018380587C2C046D8842";
    attribute INIT_24 of inst : label is "F204850214A000015493F2D3E1030843108431884020042420008000000A1EC5";
    attribute INIT_25 of inst : label is "A7AD6B110006B42529294A2140200204000A32B99E70D000E42156F08561095E";
    attribute INIT_26 of inst : label is "8D4FBAF808001B72840AAC4680FD53B0E7AF6F5BF98420000210B994A7094A14";
    attribute INIT_27 of inst : label is "0125F9004AFC300004A6000000000000000CC30500CE207902DB2C000000000C";
    attribute INIT_28 of inst : label is "00000000000000000000000000000000000000000000140A0FFFFDF800000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "C0893901166FF3AAAEFEBAEE6FA115223140844000000000020045C8C9661800";
    attribute INIT_01 of inst : label is "B99BA67F60DA392EF4F6A92F6A90F4BB699C98E779DB0C304D18B6DBFA0F09B1";
    attribute INIT_02 of inst : label is "75FDD7F7FDE864853F242ECAAC856363F2158DCFBDE3FB8FCB2CB2EE47FBF76D";
    attribute INIT_03 of inst : label is "C7F47644F973DCB5CCBBCE3328DD7DE9BFBAFF75FEFFDA19215FC901B8F9D3DF";
    attribute INIT_04 of inst : label is "6BD5FC78CE4F9C3F2B3D9ACE4FE387F57C9CFD7BF77B97F7D792F1FE5FDF5E4B";
    attribute INIT_05 of inst : label is "ACFF1FEBFFD52197E3F54865F8F8B1D58F9614B2AB55D2C296556AA4D7DFD5FC";
    attribute INIT_06 of inst : label is "CC45D61653B33C8D28FABBAF3BDAC9771AF4CD74C65FFCB3BEC870CEF6B6792C";
    attribute INIT_07 of inst : label is "FFCB2B330FD5BC57FF62C738783C6977B67B9795E489B9D6E82E54C65FFCB291";
    attribute INIT_08 of inst : label is "772EBFFFCB75D31772EBFFFCB2B338D6B1AC0783F31FF3FBFFFCB75D31FF3FBF";
    attribute INIT_09 of inst : label is "E75A985291C611BDBEA87D540A8427D73F4B72E2948E21DCFA149390B3BE3F31";
    attribute INIT_0A of inst : label is "E5737AA44AA2196208EBAC3AB579D6D7BA86C0D9E1898F269A74440000103BDC";
    attribute INIT_0B of inst : label is "5018467EB95489C03CFEDC36544CE8D4F349304C203F25F57E5CEBEE71F9C4E7";
    attribute INIT_0C of inst : label is "2D73E5A771AC4FC9B3E0E1419C02D4208100005949D5FCEABED5F75D7FD7EA23";
    attribute INIT_0D of inst : label is "1D8973E2CB25051752CB05BA2EA5960B766D8D9B67FDC366CF97D68C4CA41999";
    attribute INIT_0E of inst : label is "A42BCAAC3D2B14D65971AE48D178DD6A373097184B0C3CC75F85AD674E4C5858";
    attribute INIT_0F of inst : label is "00000000000000000000000000000000000000000000C549398CA4F815E5543D";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "BB200E06000A4000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "D9A2B20FE4ECD1518E54F3302116C88FEC8CA5CBDDE977FBEFE7DCBF0CC5784F";
    attribute INIT_13 of inst : label is "E000000000000001FC0784DBD3FC54FF153FC47637D5D85F57617DA37BD5CECE";
    attribute INIT_14 of inst : label is "524800030180DB0D900805B0D90092400030192C000041813BF77ECD16270C12";
    attribute INIT_15 of inst : label is "00000000000000000000000000000000092613060008041B6DB0000100800022";
    attribute INIT_16 of inst : label is "5015501515555051111440AAABFFA0540505AEBBBBB050400000000000000000";
    attribute INIT_17 of inst : label is "AE48DCA58A4BDAA4800580551AEEFA9106FBF106FBF106FBF106FBFEAD144005";
    attribute INIT_18 of inst : label is "A4A1884A1095CA89084538C5506A5294A4560E52D4B4210842284E5444DA0440";
    attribute INIT_19 of inst : label is "50E96068245CA5A94A5AD4A5A9084A1084A0A814E9508248A214A937394B5294";
    attribute INIT_1A of inst : label is "3F6B598E319C20FC2545AB038A108AA08ED29CE5ED6F5ED79D9C6388AE3C5126";
    attribute INIT_1B of inst : label is "2DCE0CFE1ECC331BC6D9B4426099C1084C94F9F000047A2D1461081F6B5B12BD";
    attribute INIT_1C of inst : label is "B23964D80705E1C83841D254F6A52D6B52949425084A129A4338043411C8C980";
    attribute INIT_1D of inst : label is "6309C6338E7724891324347849F3066080F6F7AFEB5ADEBFAD6738EE310227C3";
    attribute INIT_1E of inst : label is "8794A5AC4B5AE4A4A009421008F9D2448B06812A88AE006B36F465695ADEF48C";
    attribute INIT_1F of inst : label is "8DCB7586B5294A5E9484A00408501000006840A900448C12090E224502F805D1";
    attribute INIT_20 of inst : label is "800474B379303410FC21884310C431040008020A500900488D064B00758A022E";
    attribute INIT_21 of inst : label is "6100240941B686A3881708431EC6310863108631080000021000210002134153";
    attribute INIT_22 of inst : label is "5AD6BB09494A528421086054B1F34908C2A01CB5294B5294A48108DA708410A5";
    attribute INIT_23 of inst : label is "C302D0205004C3083652800528846318C621084880F044A49640A31102E92D4E";
    attribute INIT_24 of inst : label is "008532C5D93A3A7466D080C1C81714A4214A4229CB52D0CC8108C48020454906";
    attribute INIT_25 of inst : label is "9C63180100000080062108236E583AF501CC66D10810C4048D29086210862000";
    attribute INIT_26 of inst : label is "921C3380E172E49B420B12F900A81188200004012B94A58D610071842318C633";
    attribute INIT_27 of inst : label is "00047A00123C900001250000000000000008080500943A4402CF6C000000004A";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000004026000000100000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "95268D55A8924CD5D22548943B0B20D0A02D27000000000000002A2C2D280D00";
    attribute INIT_01 of inst : label is "057640919820A58998210F5210F52224963922B5AD24D6A208E60825085043CF";
    attribute INIT_02 of inst : label is "29B4A6C2B4B1496B864B41B2496CC0C1E5B30307241B606B32CB6D914B4B2080";
    attribute INIT_03 of inst : label is "B5B544D4A05991A929659CA5493736BCFB14ED29D85B4C125AE192DA6D6D7B76";
    attribute INIT_04 of inst : label is "CD0063329CA5ABAC4E7F329C90A5759959395116C2B656F173242DB15BC5CC90";
    attribute INIT_05 of inst : label is "4AAA9552A9AE435D1B6B90D746B12D48F1864896030910C912C06122A4410062";
    attribute INIT_06 of inst : label is "88CDD60C97367D8D6968CCC9735AD960889AC245C95429B6325E60DCD6B6FB2C";
    attribute INIT_07 of inst : label is "AA9B52A883E4B827CFA727BB836411CCA1A06B2489032591280810C95429B63D";
    attribute INIT_08 of inst : label is "8B5142AA9B091F28B5142AA9B52A6C6FDCDC3836432034042AA9B291F2034042";
    attribute INIT_09 of inst : label is "E58B503B6A2A226AED2B51A414AED877A9AB7A61DB516306876B28310C5D9932";
    attribute INIT_0A of inst : label is "961DDDC9B508E6EC2690BD322D77B7B7C514228019063318657242000000139C";
    attribute INIT_0B of inst : label is "CD74C36DC9E77634295FAABAFA294D0216D8251D2418E5DCB15D11EE1AC53564";
    attribute INIT_0C of inst : label is "034B0D96AE5DB2D8A5AB1DD2A1AC64D122411586B515428EA1155D7F4237FDAD";
    attribute INIT_0D of inst : label is "B794821AFCCD51E856F724B3D0ADEE4969B7B26DAC60C964AC3696EE83DA5A09";
    attribute INIT_0E of inst : label is "C686CDD500D5E20824A69B9374457A10D08004C002493CABAC14E7351C914C4C";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF02D6440CCA434366ED00";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_11 of inst : label is "3AA0006800092DB61FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "35C62767E9CAE31E53260A44C4DB76F15743AE2C313048409081324C69926352";
    attribute INIT_13 of inst : label is "600000000000000003F831242C40E71039C40E49492524A4949293C766693A3A";
    attribute INIT_14 of inst : label is "A4927924B66D24F24B66D24F24B66D37924B66D3F9361735F7EEFDEE318F8599";
    attribute INIT_15 of inst : label is "9FF9E4F3FFFF9FF9E4F3F9FF9FF9E4F209249278E097FBFE9349FCDB49A7924D";
    attribute INIT_16 of inst : label is "15155550511114414140507FFFFFAAABFFAA540505041141FFE49E79E4F3F9FF";
    attribute INIT_17 of inst : label is "2154484084216002008081415EBBBBEEAD144EAD144EAD144EAD144005501550";
    attribute INIT_18 of inst : label is "8081804A5287B8E5400C04025221084210842400020000240842495500614182";
    attribute INIT_19 of inst : label is "02148C00244810A401004010830100400084083E9D8AA8400100491204000810";
    attribute INIT_1A of inst : label is "000021000200248526E00A005082294540010000400420000210840921024422";
    attribute INIT_1B of inst : label is "12AA4004001204A409024094812042521000EDD9B36502042218C91205014242";
    attribute INIT_1C of inst : label is "20502043006114090080890810100020004010042100020085082040EAAAC085";
    attribute INIT_1D of inst : label is "8028004200800162C0813C78C084C0449020421000000850000421000000948D";
    attribute INIT_1E of inst : label is "81020082010040008520000002ECF85229021A04049415106040848500080090";
    attribute INIT_1F of inst : label is "40200240000420004000842100000084204A3CA04213E51604214C203105542A";
    attribute INIT_20 of inst : label is "183A0A313182448058008420004200042100024410A4F3E8141204B00001D025";
    attribute INIT_21 of inst : label is "2130800110908001490200010A000000210840000021000210840000000057DD";
    attribute INIT_22 of inst : label is "080106023084201004004E0020D5181001240800802000420040204A5080A129";
    attribute INIT_23 of inst : label is "0C510A250045894A101084200000C6318C631814B823A2240C28468920448420";
    attribute INIT_24 of inst : label is "180018B0306D1E3D2240293009120421080000008101004081068021DA128302";
    attribute INIT_25 of inst : label is "8001080000008484200000345418AF8FF5E44042A0AA248078006718CE718CE7";
    attribute INIT_26 of inst : label is "BD233260195D0589898009012A022000014842308100008420000214A4290A50";
    attribute INIT_27 of inst : label is "05B4020122006000122A0000000000000002A0202110021B0020008000000005";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000009048000000200000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "42845E853410066CAB52AD4A9984108AA6499B400000000002000FD151320B00";
    attribute INIT_01 of inst : label is "0576F9C37805AD499F2009F2008B2924937B7694E5249CA09A5E0125089819AF";
    attribute INIT_02 of inst : label is "A10A843A0E941B6B42DB71B6DB6ED6D48DBB5B52AD021408B2CB6DBB5B4B60C0";
    attribute INIT_03 of inst : label is "04544DD5AAC8ABAB6B6CBDAEDE33929A595082A10740E506DAD0B6DC65253732";
    attribute INIT_04 of inst : label is "186A1616BDD04023DCFD763DBA080449CB7BF3502A08D643396F810B590CE5BE";
    attribute INIT_05 of inst : label is "CB221442886C5777021B15DDC08B658065E0008150392C00102A072304D06A16";
    attribute INIT_06 of inst : label is "2A8775ACC5A5410A4F72AEEB5A5290482AB68A4A03556404A617429694A48209";
    attribute INIT_07 of inst : label is "AA8072CABD81113B3634BBD8102D3A5DC8205B7019A7655561CB9403556404A1";
    attribute INIT_08 of inst : label is "21840AAA800920021840AAA8072C45772AAD0102D0021840AAA800920021840A";
    attribute INIT_09 of inst : label is "A50AD1C2C2A4026A6420C40460888A08636A862E1615008388523100064C9800";
    attribute INIT_0A of inst : label is "9481DD8AE7B55CB6D290ED3AA351858C81E43C84A48056019472014000001294";
    attribute INIT_0B of inst : label is "03C20962FBE826AC2B41A811503BC99AE4EBADB62E5A021FB34A009032CD1565";
    attribute INIT_0C of inst : label is "6B5A4014C076E38255B2A118C80474F1A3403383B55D42AEE15D5DD542888D3B";
    attribute INIT_0D of inst : label is "13060D4420999FCAA02C002F954058004D3AC34EB001004C690025105A120C00";
    attribute INIT_0E of inst : label is "3532988CEA81C0228205E71A30D07800AC200690025941DB2D6AF7B5BDBB6465";
    attribute INIT_0F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1924D2B80114994C44EA";
    attribute INIT_10 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_11 of inst : label is "220FFEFDFEFEDF7DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_12 of inst : label is "3A1026D7018D081042A40A65FCD1A691A246302A372E4A5494A9338A499C5252";
    attribute INIT_13 of inst : label is "600000000000000000000126304488112204488919372464D49193318EDB2B2B";
    attribute INIT_14 of inst : label is "F7FA4F25B6FF64F25B6FF64F25B6FF6CF25B6FF646002245540A815187566C25";
    attribute INIT_15 of inst : label is "F24F3FF24924F24F3FF24F24F24F3FF209248049FF97FB24924FFCFE7F24F26F";
    attribute INIT_16 of inst : label is "5051111441414054015500A22288F777DDA223DDA2768DE0493CF24F3FF24F24";
    attribute INIT_17 of inst : label is "200400000100001000000FFFA505045005501005501005501005501550151555";
    attribute INIT_18 of inst : label is "00000000000458300000021012000000002100000000000000104A0000000800";
    attribute INIT_19 of inst : label is "0002020000000000000000000000000000010010C13200000002000000000000";
    attribute INIT_1A of inst : label is "8000004000002020FC180000014008004108421000000040000020083E490000";
    attribute INIT_1B of inst : label is "8000410040008000000000000000000080207CFBB76000000100090000004200";
    attribute INIT_1C of inst : label is "E2C000001082080900000802000000000000000000000004210804006A000000";
    attribute INIT_1D of inst : label is "000800000020052850A9000200000080900000000000000000000000008280AA";
    attribute INIT_1E of inst : label is "0000000000000000000000104891D24000000040208000100000040100000080";
    attribute INIT_1F of inst : label is "4000001000000000000000084000040100696A85A9F770000000811200000000";
    attribute INIT_20 of inst : label is "0A1A00000001048000000000000000000000000020A0FA18B000000108240020";
    attribute INIT_21 of inst : label is "414A10A00000101009040000000000000000000000000000000000000002D215";
    attribute INIT_22 of inst : label is "000080010842100000007172F4F0000008240000000000000000000000000000";
    attribute INIT_23 of inst : label is "000800200040000000000000000000000000000A8529F0000001004120040000";
    attribute INIT_24 of inst : label is "00412A143B670A09000006000900000000000000000000041004C0812BF80000";
    attribute INIT_25 of inst : label is "042108000000000002000024F5427E0C53600000010404820084000000000000";
    attribute INIT_26 of inst : label is "492AE014F4F80000001040000002000000842108400000000000108001004200";
    attribute INIT_27 of inst : label is "FE0E24FF87120FFFF870FFFFFFFFFFFFFFF804081E204480FC41047FFFFFFFB2";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000020D00FFFFDFC7FFFFFFF";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "468DBFF0C24B79037EFDFBF0C48C11B311347FC000000000030071EDED721901";
    attribute INIT_01 of inst : label is "30890E0C20921024498490484910849B6C94884250DB661B4D0824D8F264437A";
    attribute INIT_02 of inst : label is "1B586D6158C5A48C39246E48248F0506123C14183276B1DDC924924404228609";
    attribute INIT_03 of inst : label is "6EE5F204E3225C1484924A1021C9C841140D961B2C259169230E491B91908388";
    attribute INIT_04 of inst : label is "9ED5B8C84A0227762121894A4044EEE3A4941C89615D012C9C901B5C04B27240";
    attribute INIT_05 of inst : label is "36B3B676CEF3061336BCC184CDDC988DE1C22CB6ABC6984596D578C6B2CED5B8";
    attribute INIT_06 of inst : label is "8AD11633063661EC6080888C6388596408C0E5A4440791B6B2DB72D8C216C32F";
    attribute INIT_07 of inst : label is "555B8DA04981301326340318D8B1C3624413848666389A168CE0C6440791B6B5";
    attribute INIT_08 of inst : label is "4588ED555B969904588ED555B8DA4067008C0D8B0904588ED555BB69904588ED";
    attribute INIT_09 of inst : label is "CF1A424E72F80F971182AD30660C6328572485927397C19939C781E0392E5D90";
    attribute INIT_0A of inst : label is "62462667BD4FF7B5B8460EE767339E96CF38E71E60890024851204C000002739";
    attribute INIT_0B of inst : label is "856C4C1740BA9EFA8B2199B6DCCF264BA16D7246AF632A204C3F3650CD30C296";
    attribute INIT_0C of inst : label is "44636DE730D6BC8ABA7EE703CF04D03089049F9CC88CCC422684C4444EE8D70A";
    attribute INIT_0D of inst : label is "19084F62E261A4FB56E10DB9F6ADC21B60E4C83948C4436B0DB6D7E80E3E0C59";
    attribute INIT_0E of inst : label is "ADE7D2E7EF98C18518482241DB18810906109B884D9E42DCF1D5294E4A441051";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000071331E28026CF3E977EF";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "60800F7E000F6FBE000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "DD22D80F067691639C58F198FFB41DDC89D0618383833386670C986534C32929";
    attribute INIT_13 of inst : label is "E00000000000000000000ED9C3BC74EF1D3BC7764681D1130F646D029104CECE";
    attribute INIT_14 of inst : label is "0001B60249009B60249009B60249009B60249009BF2271F0760EC1E810FE005E";
    attribute INIT_15 of inst : label is "6DB6DB61B6DB6DB6DB61B6DB6DB6DB6009260137DF6804D96CB6D800001B6000";
    attribute INIT_16 of inst : label is "144141405401550001555000000000000055555500015541B6D86DB6DB61B6DB";
    attribute INIT_17 of inst : label is "0000000000004000000001111441450550151550151550151550151555505111";
    attribute INIT_18 of inst : label is "000000000007480001043DEE000000000000000000000000000070001043F7F0";
    attribute INIT_19 of inst : label is "43FDFDFF00000000000010000000000000000031D394002087FDC00000000200";
    attribute INIT_1A of inst : label is "00000000000000A10EB000821EBF0000000000000000004010002000254A0010";
    attribute INIT_1B of inst : label is "7000000000000000000000000000400000009429F4B001043EFFC00001000000";
    attribute INIT_1C of inst : label is "B7001043EF7DF7C00420000010000000000000000000000000002448E8002087";
    attribute INIT_1D of inst : label is "000800000000040814203E6C2087FF7C0000000000000010000000000002800F";
    attribute INIT_1E of inst : label is "00000000000000000000000002152BB800821FBFDC0000000000040100000080";
    attribute INIT_1F of inst : label is "000002000000000000000000000000200861422508536001043F7EEDF8000000";
    attribute INIT_20 of inst : label is "50A1800821FEE00010000000000000000000000000A103EDC001043EF7DBF000";
    attribute INIT_21 of inst : label is "000894200410EFEFC000000002000000000000000000000000000000000204B8";
    attribute INIT_22 of inst : label is "00000400000000000000655A84F80410F7000000000000000000000000002000";
    attribute INIT_23 of inst : label is "1FF700000000000010000000000000000000001C10020802087EFFB800000000";
    attribute INIT_24 of inst : label is "00014245992F9F361043F9FFC0000000000000000000000014A1DAD4F8500082";
    attribute INIT_25 of inst : label is "000000000000000000000036E94AFF7EB4301043FEFBE0000000000000000000";
    attribute INIT_26 of inst : label is "676FA000842800410FEFB8000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "01F1DB0078EDF000078F0000000000000007FBF7E1DFBB7F03BEFB8000000062";
    attribute INIT_28 of inst : label is "000000000000000000000000000000000000000000001F0FEFFFFDFB80000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "40841FE056DB62240A102840808010838010FF4000000000010057C7C64D1801";
    attribute INIT_01 of inst : label is "60002C4860000060090D8950D89105800110100000002C100C180000F82C0B2B";
    attribute INIT_02 of inst : label is "120848210885000810004400400E040400381010202410908000000808220C5B";
    attribute INIT_03 of inst : label is "4844A00442040838000008024081800010090212042081400204001101000300";
    attribute INIT_04 of inst : label is "9455108008422642402100080844C84280108808210802081802120808206008";
    attribute INIT_05 of inst : label is "40912224444304312410C10C4909008CE1422C12A988584582553100B0845511";
    attribute INIT_06 of inst : label is "8A531220421320A4210088882118CB24088246164006009290CF2A4846324164";
    attribute INIT_07 of inst : label is "554910242901301224340210C8A18B404416081240B000170440824006009294";
    attribute INIT_08 of inst : label is "4588E55549185904588E55549102C06500880C8A0904588E55549185904588E5";
    attribute INIT_09 of inst : label is "6B3A004E327C06160181043006006108830088027193C0B039CD90E0632A5590";
    attribute INIT_0A of inst : label is "0244006718AF9B32B42508A227339696CF21E43EE0800200811180C0000035AD";
    attribute INIT_0B of inst : label is "8420282349BB9A7E8B61332C8DE74289A1E0D866A9410A00883F24108E20A314";
    attribute INIT_0C of inst : label is "404124B2308618029C7E6703C705F06583001FB18CC44E6227CC44444C485686";
    attribute INIT_0D of inst : label is "1000CF22667194B15265049962A4CA0920E4D83908C4413E249253C1066C0C4B";
    attribute INIT_0E of inst : label is "89E33663E79CC30C30C422C1D8081318850F020780104050C0C0000008080381";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000071338E20003CF19B33E7";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "6080000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0801005E0004008210E0C020016C1B1899B22501010202040408010000080031";
    attribute INIT_13 of inst : label is "E000000000000000000008031204448111204440481101204404802080080C0C";
    attribute INIT_14 of inst : label is "180C00DB0180C00DB0180C00DB0180C00DB0180C00C871E02204408109FA040F";
    attribute INIT_15 of inst : label is "0000000C00000000000C00000000000C09276580000804020100000180C00DB0";
    attribute INIT_16 of inst : label is "40540155000155555400000000000000000000005555554000030000000C0000";
    attribute INIT_17 of inst : label is "0000000020000000042005050140411555505555505555505555505111144141";
    attribute INIT_18 of inst : label is "4001000000068D00000000000008421084108040100400000200000000000000";
    attribute INIT_19 of inst : label is "000000000000000000000000010000000000002881A000000000000000000000";
    attribute INIT_1A of inst : label is "4000002000000000040000000000000000002108000000000000000000000000";
    attribute INIT_1B of inst : label is "000000002010042008020084010002104000E902000000000000000000000000";
    attribute INIT_1C of inst : label is "60800000000000000000000100000000000000000000000210003B0284000000";
    attribute INIT_1D of inst : label is "0000000000100122408142840000000000000000000000000000000000001760";
    attribute INIT_1E of inst : label is "0000000100001000000000007684081000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "00000008000000000000010422008000004912040A1420000000000000000000";
    attribute INIT_20 of inst : label is "D5A10000000000000000000000000000000000020005D8182000000000000000";
    attribute INIT_21 of inst : label is "004810200000000000000000000000000000000000000000000000000000157A";
    attribute INIT_22 of inst : label is "0000002084210800000049020508000000000000000000000020000100000084";
    attribute INIT_23 of inst : label is "000000000000000000421084210884210842104001D3A0000000000000000000";
    attribute INIT_24 of inst : label is "000048903070A142000000000000108421084200000000000408800100000000";
    attribute INIT_25 of inst : label is "000000000840000001000020C10283D7A7400000000000000000000000000000";
    attribute INIT_26 of inst : label is "66E7800025000000000000000000000000000080000000200000004210800000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000062";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000FFFFDF800000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
