-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FD7CF75BDF7F7BEBDF534F7F53DBDF7DFDEFEF7F55EDD6F7FAA08A2088834699";
    attribute INIT_01 of inst : label is "7BEBDF53D5FDF34BDF7FF5FFAFFD55DF3B7DD2FFDBDF5EFAF7D4D3F74BDF7F7E";
    attribute INIT_02 of inst : label is "CD7DBDF5EBD4F3B3B34F6F6F7D7BEBDF535FCD2F7DFFD7FEBFF575ECD2F7DFFD";
    attribute INIT_03 of inst : label is "34FDD2FF7FD7BEBDF534ECFDD2F7DBF7EFD7CD3CF6F7D7AF53CF3CD2F7D7EFD7";
    attribute INIT_04 of inst : label is "FD7FEBFF5573DED4BFF6FFF7FFBFFD34FCD6FFDF5EBD5F7CF3DD2F7FD7BEBDF5";
    attribute INIT_05 of inst : label is "6FEF7D7BEBDF535FCD2F7FF7D7BFBDFD74FD5BDFFDF5EFAF7D4F75B7DF52F7DF";
    attribute INIT_06 of inst : label is "FEBFF574EDF74BFF6FDFBF4D7DBDFDEBD5D77CBDFDFBF5F35F6FFF7EFD7CD3CF";
    attribute INIT_07 of inst : label is "FDFBF4ECF7F75F6FFDF5EFAF7D4F75B7B34BDF7FF5FFAFFD55CF3F572FFFFFD7";
    attribute INIT_08 of inst : label is "F35B3CEDBDFDEBD5D7CF6FFFF5FFAFFD54EDECF3CD2F7DF5FBF4F3B3CD3CF6FE";
    attribute INIT_09 of inst : label is "3DF56FFDDD7FEBFF57CF3D5CF7CF52FFDF7D7BFBDFD57B573B6F7FBF7EFD7CED";
    attribute INIT_0A of inst : label is "3B7B53F2F7DF5FFAFFD55CF34BFF6F7D7BEBDF535CFD4BDF7DFDEFEF7F55DF7F";
    attribute INIT_0B of inst : label is "F575B3CF3D4BFF6F7D7BEBDF57CD73B35CBDF7FF5FFAFFD55CECF34BDF7D7EFD";
    attribute INIT_0C of inst : label is "77CF52FFFF7D7FFBFFD7CF57B35DF6F7DDF7FEBFF5573B7F56CF2FFFFFD7FEBF";
    attribute INIT_0D of inst : label is "F5FFAFFD55F3CFDF572FFFFF5FFAFFD5D73CF7DDECD2FFDBDF5EFAF7D4D7DF77";
    attribute INIT_0E of inst : label is "F7FFDFBF4F3DDF77735BFBFFDFFEFFF4D7D5BDFFDF5FFAFFD5D6CF7F7DD2FFFF";
    attribute INIT_0F of inst : label is "6F6F7D7BEBDF535DCF73B777D4B77D7AF556CFCF76FFDFDEFEF7F5F75CFD5F76";
    attribute INIT_10 of inst : label is "EFDFBF4ECF7F75F6F7D7AF57F3CF7F52F7D7EFD7DDED5F76F7F7AF57DDD3DDF7";
    attribute INIT_11 of inst : label is "F53DF7CD2F7F7EFD7F3B73DF7756DD7AF57CF3D377CF52F7D7EFD7CCF7573B6F";
    attribute INIT_12 of inst : label is "F7B3CEDED4BDFFDF5FFEFFF4D3B3B756F7FF7D7FEBFF55773B7773B52FFDBD7A";
    attribute INIT_13 of inst : label is "53B577D4ECBFFFD7AF57DCF735DCF776F6FDFBF5F73DD5F73CBDF7D7FEBFF553";
    attribute INIT_14 of inst : label is "AAAA845551555440000BFFDFFEFFF4D3B73F3D5BDF7F7AF57D4FDBFFFD7FEBFF";
    attribute INIT_15 of inst : label is "111111111111111111111111111111111111111111111111110111111108AAAA";
    attribute INIT_16 of inst : label is "25296BDEF7D8E6218E63D695B5ED6DC8631EB5AD2F7BE5B4B9B2151111111111";
    attribute INIT_17 of inst : label is "C4294838C6309CE5B1CC7310C6A56B6BDADB98C729487356B4BDAF7D8E621486";
    attribute INIT_18 of inst : label is "B5B631CE4290E6A56B7BDEFB9884318E7A56B7BDEDB9885398718C2739CF739C";
    attribute INIT_19 of inst : label is "F6BDEDB98E6398E63D694BDEF7DCC7318A639EF4A5296BE85218E6398B4AD2D7";
    attribute INIT_1A of inst : label is "42308CE52DCE6318E639EB4A5696BEC73988531CD4AD2F6BDF6318C5298E6A52";
    attribute INIT_1B of inst : label is "521EB5AD2F7B6E6398C531CF7A5294B5F731CC721CC38C63294E7B98E639CC61";
    attribute INIT_1C of inst : label is "9990A273998CC8403C88C5281C05901EFB42B98E6398E63D694BDEF7DCE7310A";
    attribute INIT_1D of inst : label is "8CA05038CC0201CCE6722144C623194826399CCA4131CCE50289CE6472890E73";
    attribute INIT_1E of inst : label is "45129CC4720904C73140A007399C884131CC8E44218E4728144E7339900A7311";
    attribute INIT_1F of inst : label is "738F33C4F9CE318CE33E3398E633C738CE38CA71C651C6719CEA18A975D7FCCC";
    attribute INIT_20 of inst : label is "650CA500CA96427BED28028802799CF399E7C7319C6718E78C638CE71CE318C6";
    attribute INIT_21 of inst : label is "208A110659401204B2804594032942194A01943208B204A01167290022864190";
    attribute INIT_22 of inst : label is "4B6C97F5DFD6082B0882208A280240842294211065284220CA50804194A10883";
    attribute INIT_23 of inst : label is "700700700700700700E1A43D7555FFD4F752AAAAAA44E28595CBBAFFA24924B6";
    attribute INIT_24 of inst : label is "66556D365071669204010C431040310C4100C431040310C41700700700700700";
    attribute INIT_25 of inst : label is "A8F6169EEDAAF618A8336777726167537577C324628430624724124720325661";
    attribute INIT_26 of inst : label is "0B84B3A8493AA1D8FADBBEA9D8E281BFE7EAE638AE6382B40C0B5080B48C0ACC";
    attribute INIT_27 of inst : label is "69DA969DE0A6C865B298E1B79D7BB618A9B68C3B87D79FE998F6DB9EC8D0B40D";
    attribute INIT_28 of inst : label is "4872902FDE5BF796FDE585E938D2F3BD7F9FD2D3B56D3FC2B0BC6979DEB7CDE9";
    attribute INIT_29 of inst : label is "24820924820924820924820924100400A242A653A53C0429485290A5211CA439";
    attribute INIT_2A of inst : label is "9E09E0DE0EE0EE0EE0EE0EE10040083684210825029249248209248209248209";
    attribute INIT_2B of inst : label is "761F8761D8761D87E1D87E1F87E081D8053C0F60EE0EE0DE0EE0EE0EE0EE09E0";
    attribute INIT_2C of inst : label is "210052108521085A1084A10852108521085210852100C0210461D87E1D87E1D8";
    attribute INIT_2D of inst : label is "9CC731C100212082082080069A69A69A0020820820EBAEBA638E3801CF3CF3CF";
    attribute INIT_2E of inst : label is "605041E0683B0EC3B0EC1E0404801811C16C11C11C0482A5210A5210A5080200";
    attribute INIT_2F of inst : label is "14050180701807018040280780380380380E80D80380D80E820301C1185E1184";
    attribute INIT_30 of inst : label is "3903403402C00C04D05505D0490810000300C0100C0100C0100C0100C0101060";
    attribute INIT_31 of inst : label is "061A697AA474D8083A0C0280C030148421285210741805018060350942509410";
    attribute INIT_32 of inst : label is "804A89414867A333DA4F25333331C809BCE4CAFF4333D99FF2EC970BA96FEFE1";
    attribute INIT_33 of inst : label is "EAB26B11E3E7FB0EDF2B0422C211410810810E0C0001932F407825333331CCE5";
    attribute INIT_34 of inst : label is "A6DF17EB7973FB3FA60A24133270F2D667256E11DD60920BDDE45DF6AB9EA3AA";
    attribute INIT_35 of inst : label is "BCEF36799F7BBEAEF2231853C89F956E4C08A0C354EA908651F5CEFF387C7F07";
    attribute INIT_36 of inst : label is "F7D3ADB2F08DD2DCABFAE5D7860F2AD6C3D00DE956482186CFF9604D45AEC026";
    attribute INIT_37 of inst : label is "FE2C53CC9F6DC17C27A8DC773C1AFB448122938A9E5267ACECF1BAF875A04F8E";
    attribute INIT_38 of inst : label is "14D43DC4803430190960000422002012BB7DDE9FFDCBFD1DFFF37FFFFFFF7FE5";
    attribute INIT_39 of inst : label is "210A2650881912250000402000D14406B4FB5BC0FAFFFDFF7EFE6FFFF1FFDFEF";
    attribute INIT_3A of inst : label is "C14461E07058020081C2405C52A41802D6F5EAFD9D6FEFD69E68FB7AEB7A97F1";
    attribute INIT_3B of inst : label is "2E2C02200C145030570D2C2020165401A3327F77BE7FF1A2B78B0B6F9FF4FEFF";
    attribute INIT_3C of inst : label is "C80209038D03CCE000880080005A0104FF778FBADDCFA7CA7FFBFF979F37FC7F";
    attribute INIT_3D of inst : label is "080256080009D86400A20020700C8242FE6DDFDDB79FF3FFFFDDFDFFFD7DFFFF";
    attribute INIT_3E of inst : label is "29512D9C06001C0CA492B80509BA86FB5FBEFE8EE39BD8DF9AFD93F45DAF7FAF";
    attribute INIT_3F of inst : label is "8C8841C182EF011A0BE013104C2A457525B7F9279F9167E5E51AEADEFFF6BFF7";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "F95D71D3EF3E7DE3EF11D75D71D3EFBEF1E78F3C5D7570F3CFF9E3C75B072CB2";
    attribute INIT_01 of inst : label is "7DF3EF91DD7571D3CFBEF9F7CFBE5DD7195C74FBEBCF9E7CF3E475D5D3CFBE7C";
    attribute INIT_02 of inst : label is "D75C3EF9F3E575D5D5D74FAFBC7DE3EF11D7470F3EF3E79F3CF95D6574FBEFBE";
    attribute INIT_03 of inst : label is "5C7470FF3FE79F3CF91C757474F3EBE7CF95C71D74F3E7CF91D71C74FBE78F15";
    attribute INIT_04 of inst : label is "3E79E3CF1775D65C3CF2F3C79E3CF11D6570F3EF9F3E575D75D74F3FE79E3CF1";
    attribute INIT_05 of inst : label is "4FAF3E79F3CF91D7574F3CFBE7DE3EF15D75C3CF3EF9E7CF3E475D95C774FBEF";
    attribute INIT_06 of inst : label is "9E3CF11D6575C3CF2F9F3E471C3EF9F3E4771D3CF1E3C575C74F3E7CF91D75C7";
    attribute INIT_07 of inst : label is "F1E3C47575D5D70FBEF9F7CFBE575DD5D5D3CF3CF9E78F3C5DD71D774FBCFBC7";
    attribute INIT_08 of inst : label is "75DD5D753CF1F3E471C74FBEF9F7CFBE5D757575C74F3EF9E3C475D5D75D74F2";
    attribute INIT_09 of inst : label is "5D774F3CEE79F3CF95D75DDD75D774F3EFBE79E3CF1759775D4F3CBC78F15D75";
    attribute INIT_0A of inst : label is "5D5D71D4F3CF1E78F3C5DD71C3CF2F3C79E3CF15DC65C3CF3CF9F7CFBE5DC75D";
    attribute INIT_0B of inst : label is "F91D95D75DD3EFAF3E79F3CF95C775D5DC3EF3EF9F7CFBE5DC7571D3CFBE78F1";
    attribute INIT_0C of inst : label is "75D774F3CFBE79E3CF15D77595DD74FBCEC7DF3EF9775D1D77570FBEFBE7DF3E";
    attribute INIT_0D of inst : label is "F9E78F3C5D75D75D774FFBCF9E7CF3E5775D775D7574F3EBEF9F7CFBE575D777";
    attribute INIT_0E of inst : label is "F3EF9F3E471DD77775D3EBEF1F78FBC5765C3EFBEF9E7CF3E577575D1D74FFBC";
    attribute INIT_0F of inst : label is "4FAFBE7DF3EF95DDD775D775DD3BBE7CF977464774F3CF9E7CF3E575DD75D770";
    attribute INIT_10 of inst : label is "2F1E3C47575D5D70FBE7CF95D5C75D74FBE78F11DD75D774F3C7CF95DD75DDD7";
    attribute INIT_11 of inst : label is "F11D75D70F3E7CF95D5D75DD7774EE7CF95D75D175D774FBE78F11D577775D4F";
    attribute INIT_12 of inst : label is "D5D5D7575D3EFBCF9F7CFBE475D5D774FBEF3E7DF3EF97771D7771D74FBEBC78";
    attribute INIT_13 of inst : label is "95D775DD753EFBE7CF95DD775DDD7774FAF9F3E5775DDC775C3EF3E7DF3EF975";
    attribute INIT_14 of inst : label is "5555541554540500000BCF9E7CF3E571D75D5DD3EFBE7CF95DD743EFBE7DF3EF";
    attribute INIT_15 of inst : label is "1111111111111111111111111111111111111111111111111101111111375555";
    attribute INIT_16 of inst : label is "10C610040058C73908431CC6214A45CE52084210800027EB18723CD111111111";
    attribute INIT_17 of inst : label is "C739CC6318E72108B9CC7318A310C410002B1CC7398C5318C62908458C6398C4";
    attribute INIT_18 of inst : label is "0817318E73988631CC42148B98C729083108400842B18E6294C631885291739C";
    attribute INIT_19 of inst : label is "842148B98C7398A4398E6290855CC6398C4218C631CE522C7310842144210820";
    attribute INIT_1A of inst : label is "88431802058E631484298C6318E522E7398E6214E639884211731CC739486398";
    attribute INIT_1B of inst : label is "73084218C0002E631CC6210C6318E7291631CC731486318C42108B18C7318E51";
    attribute INIT_1C of inst : label is "0898C46201404E633440863918BF2EF04504B98C7398A4398E6290855CE731CE";
    attribute INIT_1D of inst : label is "40C462340F33118880503188C412818C6728100C6331008623118A2243118E42";
    attribute INIT_1E of inst : label is "062318A0439988E4298CC44620100C633904080639880439988C41281C8C7281";
    attribute INIT_1F of inst : label is "779F73DCFBCEF3BCEF3EF3B9EE77CF79DE7BCAF3DE57CEF3BCE21289D7DDD008";
    attribute INIT_20 of inst : label is "85B0A60B0979F984544400A002F9BCF79BE7DF379DE779EF9DE7BCEF3DE779DE";
    attribute INIT_21 of inst : label is "2B0B21585B8260B8330585B8242B83614C161642B0B704C1616C2982C2D85215";
    attribute INIT_22 of inst : label is "9001257F5DF5DF5DB0A42B0B704C170642B8361485706C290AE0DC1215C1B0A4";
    attribute INIT_23 of inst : label is "28028028028028028010BEC42BBB1115B946BBAFFADB07FF15BFAEBEE4800000";
    attribute INIT_24 of inst : label is "CA2292EB2186FA65840101C070180701C0601C070180701C1280280280280280";
    attribute INIT_25 of inst : label is "F28125291AD1896B3832C9AF95DFBE75D7BFE7968B2692CB2282EA2686DA6282";
    attribute INIT_26 of inst : label is "624004348653C0063484434C272C418C39DBDBDFBDBDB389EF1896B399EB189E";
    attribute INIT_27 of inst : label is "1018A1010080524938E04834824834800F3C104806988535A94A52D680042080";
    attribute INIT_28 of inst : label is "91B52024FBE93EFA4FBE858E30880730C41108E600CE61028109C86080A43908";
    attribute INIT_29 of inst : label is "8A28A38E38E28A28A38E38E28A100400EDF75B2430C904EB19D633AC616D48DA";
    attribute INIT_2A of inst : label is "6E06E02E00E01E00E00E00E10842082A8421082B0238E38E38E28A28A38E38E2";
    attribute INIT_2B of inst : label is "060580601806038160181605816080981F6402601E00E02E00E01E01E00E06E0";
    attribute INIT_2C of inst : label is "210016038160780E0380E03816038160381603816100C0210060181603816018";
    attribute INIT_2D of inst : label is "58F7B5A10020268A68A68825105105120A48248248840040B4C34C8292092092";
    attribute INIT_2E of inst : label is "A040408000010340100408040400700340340340340402108C6318421090E729";
    attribute INIT_2F of inst : label is "08020000200002000040F80C80D80D80D80480180D801804820E0300280A0280";
    attribute INIT_30 of inst : label is "1304F04705707703702F03303F08100201800010000100001000010000101000";
    attribute INIT_31 of inst : label is "ED3D923CDAA961081611846178460781603816102C2308C2709C0B06C1B06C10";
    attribute INIT_32 of inst : label is "1964C98B037E49818E0621AAAAA3A7B9AD4AF52A89818C0CD2404671C82C4443";
    attribute INIT_33 of inst : label is "133022916687D487905477563B8D3DC7DD7DC7250002DBF89DFAA1AAAAA3AFCA";
    attribute INIT_34 of inst : label is "DBBDFEB08BF0B78D662D7F3F5EFFF2DA424080070718022051B14180414E7D05";
    attribute INIT_35 of inst : label is "F7BFFFFDFEBEB6DEB5383B2BDF57FC7B15021800585182A0066C44C992000084";
    attribute INIT_36 of inst : label is "8420A14A05A3905444244508210045907BFF9F7EDCDCDCD87FF7FFFEC75FB5BF";
    attribute INIT_37 of inst : label is "0D4809058000330B04C0221082188271ABAFFF6F53D6AF55B9FFA7A77B36FFFB";
    attribute INIT_38 of inst : label is "47084405A5856108320100DC08290091D9D3FFDFBD505FA5FFBAF7FF4F5FEFFF";
    attribute INIT_39 of inst : label is "65000C310C83907000810105321BC880FCEA5ED79AD7C7EFD6A8FFA8BFBAFFFD";
    attribute INIT_3A of inst : label is "5FDAFABFFFE7FDF8D7FD609E9FA71D970AA009004196421C6023388832F80701";
    attribute INIT_3B of inst : label is "93743BFFB3FBF63D7C75F17F6BCB1FD30082227288008842044D020CA0059821";
    attribute INIT_3C of inst : label is "56C50CA8C6718012A091107D02003E0CE7CDBB6F6DF3D72D8A97FE1B558DFFFB";
    attribute INIT_3D of inst : label is "2750400720E29A2E20AC124251C140061F7F6FADFBF9D4DD9FFBFFFDAF8D23C6";
    attribute INIT_3E of inst : label is "FBEBBFAD7FD99FFF3BBBF7FFF73A32B3051009A24004112105885F0880449B80";
    attribute INIT_3F of inst : label is "5F9BF3FDEACFBFFF7B7DF5DBD4B6CFBE25960040B82A3441434046081CDC0D01";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "B15C7542EBAC5D62EB15471D55C2CBACB975CBAE546554BAE001FD43E55270E1";
    attribute INIT_01 of inst : label is "5D72EB95D4647552EBACB1758BAC55C75D1D50BACACB965CB2E555D152CB2C58";
    attribute INIT_02 of inst : label is "D55C2CB972E4719191470BAB2C5962CB1146550BACBAC5D62EB1157450B2EB2C";
    attribute INIT_03 of inst : label is "557554BB2EC5D62EB155646450BACAE5CB91C55D70B2E5CB95C71D54B2E58B11";
    attribute INIT_04 of inst : label is "AC5962CB1571C6542CB2BAC5D62EB1557450BAEB162C471C71C50B2EC5972CB9";
    attribute INIT_05 of inst : label is "0B2B2C5962CB1146450BACBAC5D62EB1157542EB2EB1658B2C5715D1D750BACB";
    attribute INIT_06 of inst : label is "D72EB914747152EBAB972E555C2EB972E5575D2EB162C475474BAC58B15C51D7";
    attribute INIT_07 of inst : label is "B162C5647191474BAEB1758BAC5715959142CBACB175CBAE55C759570BAEBAE5";
    attribute INIT_08 of inst : label is "71591C642EB962C455D74BAEB1758BAC54646471C50B2EB162C47191C51C70B2";
    attribute INIT_09 of inst : label is "1C750B2E8C5D62EB11C71D5C71C750B2EBAC5962CB151D57190B2CAE5CB91C64";
    attribute INIT_0A of inst : label is "59195594BACB975CBAE55C7152EBABAC5D62EB155D7542EBAEB1758BAC55D719";
    attribute INIT_0B of inst : label is "B115D1C71D42EB2BAE5D72EB91D571955D2EBACB1758BAC55D647542EB2C5CB9";
    attribute INIT_0C of inst : label is "71C750BACBAC5962CB11C751D15C70BAC8C5D62EB157195956474BAEBAC5D62E";
    attribute INIT_0D of inst : label is "B1658B2C5471C659574BBAEB1758BAC4571C765C6450BACAEB1758BAC451C777";
    attribute INIT_0E of inst : label is "B2EB162C575DC7777142CAEB1758BAC457542EBAEB1758BAC45647195C50BBAE";
    attribute INIT_0F of inst : label is "4B2BAC5D62EB115DC7719771D423AC58B156575774BACB1658B2C4715C654774";
    attribute INIT_10 of inst : label is "2B162C5647191474BAC58B1591D71950B2C5CB95DC655770BAE58B11DC51DD97";
    attribute INIT_11 of inst : label is "B15C75C50BAC58B1191971D977508C58B11C71D571C750BAC58B15C57757190B";
    attribute INIT_12 of inst : label is "9191C646542EB2EB165CB2E451919754BACBAC5D62EB1577597775950BACAC58";
    attribute INIT_13 of inst : label is "159571D4652CB2C5CB91DC7715DC7770BAB972E4771DD5771D2CBAC5D62EB151";
    attribute INIT_14 of inst : label is "FFFFF66777677640000AEB1758BAC45597591D42CB2C5CB91D5652CBAC5D62EB";
    attribute INIT_15 of inst : label is "55555555555555555555555555555555555555555555555555455555557FFFFF";
    attribute INIT_16 of inst : label is "6318C6B18D5485210A4210852148454A5210842108529C50196738D555555555";
    attribute INIT_17 of inst : label is "A5214A4214A42108A9085290AD6318D6358A1484290A5421094A52850A4294A5";
    attribute INIT_18 of inst : label is "6315214A5294A5210A52908A14A4290A5290A42148A948521508421084215214";
    attribute INIT_19 of inst : label is "84210AA10A4294A5635AC6B58C5085214A429084214A42284290A4215AC6B18C";
    attribute INIT_1A of inst : label is "25294250850A5294A42B18C631AD62A42948421484210842154214A5210A5290";
    attribute INIT_1B of inst : label is "529085290842284290A521508421294214214A42948D6B18C6B18A10A4210A54";
    attribute INIT_1C of inst : label is "00108042090408403400852010ABAFBEAFEBA10A4294A5214A42948454852948";
    attribute INIT_1D of inst : label is "00A050300D120100A0512900850281080520144A402944840201082042094A42";
    attribute INIT_1E of inst : label is "24029480528144842904800420900840210048042948042810484028940A4201";
    attribute INIT_1F of inst : label is "BDCF9DF67CF7B9CF7B9F3DECF3BDE79EF73CF3B9E79DE73DEE6A3A0B7777D008";
    attribute INIT_20 of inst : label is "056098040801501404040200033EEE79EEF3E7DDCE7BDCF3EF73CF7B9E7BDCE7";
    attribute INIT_21 of inst : label is "240AC12056018240AC020560182402C13008158242AC03008158260102B04C12";
    attribute INIT_22 of inst : label is "924924280288808B6098240AC030480582402C13048058260900B04C12016098";
    attribute INIT_23 of inst : label is "D41D41D41D41D41D4100FAFBD4141545FEF85041449B34434E81444510124924";
    attribute INIT_24 of inst : label is "2D3CEBAE36DB0C3C84210F03C0F43C0F03D0F03C0F43C0F01D41D41D41D41D41";
    attribute INIT_25 of inst : label is "BAD6B9EE739AD6B1E82AA2CAA0820828A2EBB2D31DF9F7DF75C77C79E79E74D3";
    attribute INIT_26 of inst : label is "FFED7BDF5FDFE918C719CE6158C7814A5A9084214A5AD8D631EE739AD6B1EE77";
    attribute INIT_27 of inst : label is "0110E129C08821820C134A2872C728A3010CB0C704856A5090850D6A6579DF5B";
    attribute INIT_28 of inst : label is "7CDEF83B0496C125B049058800042111025094400046708246310E51804709C6";
    attribute INIT_29 of inst : label is "38E38F3CF3CF3CF3CE38E38E38108420B08980B8A888840C6018C0318137BE6F";
    attribute INIT_2A of inst : label is "0408403402C01402C0AC0AC10842080C0401002B00F3CF3CF3CF3CF3CE38E38E";
    attribute INIT_2B of inst : label is "5C058140505403014070141505408098098602601402C0B402C01409402E0040";
    attribute INIT_2C of inst : label is "41000601806038060181E01806018060180601806100C0318060701413014070";
    attribute INIT_2D of inst : label is "D084296108200830C208300E3CF38E3C028B2CA28B1C61871C61870082492082";
    attribute INIT_2E of inst : label is "611840A0BC0701C0701C2B0401813C01C01C01C01C11C2C6318C639CE7000010";
    attribute INIT_2F of inst : label is "0C03004020080200404048008078008078048058008058048205046018060180";
    attribute INIT_30 of inst : label is "1200A01601A00201E00700201308000000802000020000200002000020001020";
    attribute INIT_31 of inst : label is "6F06DB4F6C6D880814070140300C070160700610280E028060180E00C0200C10";
    attribute INIT_32 of inst : label is "1180FB8202081BC89C02109999918B115718142203C89C0409054152F0055443";
    attribute INIT_33 of inst : label is "049A00E71CD9100F60C48CCC06422322332326422A28005418FBD09999918158";
    attribute INIT_34 of inst : label is "7075A7FDF5DFE278BF7F98CC3D765FBB2060A782C044B10459AB688319444445";
    attribute INIT_35 of inst : label is "73EFFEEFB3F7C73EA674BCB7BEADF5B26AECA0060C4406151503424A408502AA";
    attribute INIT_36 of inst : label is "047740E2618582A161183068500261ACE986B98A69DB1F79C6BFF274FCFDB6FD";
    attribute INIT_37 of inst : label is "A01D690558990119C0450905404B9205A6BB63FB5ADF1FBAEFFBECB4FDCEF279";
    attribute INIT_38 of inst : label is "00E5488E20268001B410080474160090CFEDFAB96BA6F9BBF8CEDF5EFEBFFF2F";
    attribute INIT_39 of inst : label is "01481313C3154A00558CC602440000109CF8AF93FDBDD2DCBF27FD42FDEBF927";
    attribute INIT_3A of inst : label is "CF8FFDCEECA4FFDFEE6D7F5C38FF5EAD40010C02438088118612250490801287";
    attribute INIT_3B of inst : label is "BFFEF9FFCADAB6F6C3D2AE37F9EE7BBA44031006912104E6006D232581C936C3";
    attribute INIT_3C of inst : label is "E0580302100100E4204800490A02A842FF9E9AD733FDEF76954E6DE5DAFFE77E";
    attribute INIT_3D of inst : label is "80112125308000AA834202201285A20043F1E682DEFB6D47FFC6CFA7F7DFF55F";
    attribute INIT_3E of inst : label is "FFFFE1F1EFEB7F675BD2D3FFFFDEBFFB10529402180D110546A4800349001904";
    attribute INIT_3F of inst : label is "D7DFFF6EF7EFDFB7F6EFE7FCBA6975FA055044490452340118A52C3030493011";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "508A2CA165142CB16588A288A8A1459450A285142B2228514551BAF90457FF00";
    attribute INIT_01 of inst : label is "2CA16508AA2228A1459450A285142AA2888A285149450A2851422888A1451428";
    attribute INIT_02 of inst : label is "A28B1650A143288888A28525962CB1658CA222C51651428A14508A2328516514";
    attribute INIT_03 of inst : label is "8A22285515428A14508A222328514962C588B28A2859428508A2CA2859428508";
    attribute INIT_04 of inst : label is "1428B1458AA8A32B145A5962CB16588A222C59450A1422CA28A28515428A1450";
    attribute INIT_05 of inst : label is "85A51428A1450CA23285165142CB16588A22B1459450A28514228A88A2A85165";
    attribute INIT_06 of inst : label is "CA1650CA2228A165258B16328B1458A1422ACA1450A14228B285162C58CA28A2";
    attribute INIT_07 of inst : label is "58B162222888A2851450B28594228A8888A1651650B2C5962AA288AAC5145142";
    attribute INIT_08 of inst : label is "28A88A221458A14328A2851650A285142A222228B2851450B1632888A28A285A";
    attribute INIT_09 of inst : label is "8A2A8596442CA16508A28AAA28A2A859451428B1458AC8AA888516962C588A22";
    attribute INIT_0A of inst : label is "8888A88859650A285142AB2CA14525962CB16588AA22B1459450A285142AA288";
    attribute INIT_0B of inst : label is "50CA88A28AA16525942CA16508A2A888AA1459450A285142AA2328A165942C58";
    attribute INIT_0C of inst : label is "A8A2A85165142CB16588A2A888AA28516462CB1658AA8888AA2285145142CA16";
    attribute INIT_0D of inst : label is "50A2C5162A28A228AA8559450A2851422A8A2A2A22285149450A28514228A2AA";
    attribute INIT_0E of inst : label is "59450A14228AA2AAA8A149458A2C51632A2B1451450A2851422A22888A285594";
    attribute INIT_0F of inst : label is "85251428A14508AAA2A88AA8AA11142C58AA2222A851658B2C596228AA22A2A8";
    attribute INIT_10 of inst : label is "A58B162222888A285142850888A288A85942C588AA22A2A851628508AA28AA8A";
    attribute INIT_11 of inst : label is "588A28A2C51428508888A8A8AAA84428508A28A8A8A2A85142C588A22AAA8885";
    attribute INIT_12 of inst : label is "8888A2222A1459450B28594328888AA851651428A1450AAA88AAA88A8514962C";
    attribute INIT_13 of inst : label is "888AA8AA22145162C588AA2A8AAA2AA85A58B1622A8AAA2A8A1659428A1450A8";
    attribute INIT_14 of inst : label is "0000292C382C2C000009450A285142288A888AA1451428508AA231451628B145";
    attribute INIT_15 of inst : label is "AABBABBAABBBBBAAABBABAAAABABBABAAABBBBBABAABAAAABBBABBBAAA800000";
    attribute INIT_16 of inst : label is "425284A108508529485631AD635AC50A5284200842003FFFE288C66AABAABBAB";
    attribute INIT_17 of inst : label is "84210884A1294212A108529480084200002A9085294844A5084A108548421084";
    attribute INIT_18 of inst : label is "0014214842108C6358C6318A148421481004200042A148521421004210015290";
    attribute INIT_19 of inst : label is "210800A10A5210846B18C6B1AD508529085200000000002A5214842900000420";
    attribute INIT_1A of inst : label is "10852948550A52148428020004200A84294852918D6B5AC6B14214A421480080";
    attribute INIT_1B of inst : label is "420020084000A842948429108421084214214A5290A94A5094250A9484214842";
    attribute INIT_1C of inst : label is "AA34A8D623051A413540856291FBBEFAEAFBA10A5210844A1084A12954A42108";
    attribute INIT_1D of inst : label is "418A44301C02011188D42151A412035A2C223118C16111AD52A358AA46AB0AC6";
    attribute INIT_1E of inst : label is "0546B582568B01856154A8046A350A5161510AA42908A46A9518D56A3008D601";
    attribute INIT_1F of inst : label is "38EF98E33C633CC671DF38CE7118F78CE79C671DE718F339C72038837F5DF51A";
    attribute INIT_20 of inst : label is "0B6358F61401501551500000033C4739CC79E389E6719EF3C63BCE73DE739EE3";
    attribute INIT_21 of inst : label is "5636C2B1B63D8763EC7B0B63D8561EC2B1EC2D85616C7B1EC6D8D63D8DB1AC6B";
    attribute INIT_22 of inst : label is "000000820220A8A961585616C3B0EC7D8D63EC2B0AC3D856358FB1EC2B1F6158";
    attribute INIT_23 of inst : label is "08008008008008008054FBEFEBBBFBFE55414111040000000001504040000000";
    attribute INIT_24 of inst : label is "104114704924934904210280A0280A0280A0280A0280A0281080080080080080";
    attribute INIT_25 of inst : label is "810842118C25294E502210410E38E38E38C20008600000410C20C20820E20104";
    attribute INIT_26 of inst : label is "211AC6212862062108663096A53961010846318C631880008401004631884318";
    attribute INIT_27 of inst : label is "7284463100B8E20C30A28F3C11433CF2CA30E18204A4200A4621A86302020024";
    attribute INIT_28 of inst : label is "23004020208008200208040443188429C2309CA529884002420084021CE5194E";
    attribute INIT_29 of inst : label is "14514410410410410410410410100400A490C72CB24305C233846708C1C01180";
    attribute INIT_2A of inst : label is "9E01E0360AE03E0AE02E02E10040080D04010023005145145145145145145145";
    attribute INIT_2B of inst : label is "0E01816158160784603846018060803809BC00E03E0AE03602E0BE03E02E01E0";
    attribute INIT_2C of inst : label is "C1001A0681A0681A0681A0681A0681A0681A0681A100C0310060384607806138";
    attribute INIT_2D of inst : label is "0A4210810820B8E38F3CF00C30C34D34038E38F3CF0830C30830C30020820C30";
    attribute INIT_2E of inst : label is "C07840201C0300C02008030407806C06C06C06806807C2421084210842358C63";
    attribute INIT_2F of inst : label is "0E0380208C2B008020404817C12C13C12C01815C13C05801820501E0781E0701";
    attribute INIT_30 of inst : label is "0701F01701B00F00B01301F013081C178461185E1185E1185E1185E1185E1028";
    attribute INIT_31 of inst : label is "E912CB6A2C8D8808020280A008020481A0681A1004050140D0340D0140501410";
    attribute INIT_32 of inst : label is "01ACA342050A5300980203333331A874AC4E117DC3009805147C0D7AA6FFBFBA";
    attribute INIT_33 of inst : label is "7DB152F94FB4BA9A12D461D130CC98678778676B00082840A3F903333331A112";
    attribute INIT_34 of inst : label is "550F9DCF3E5A3745A6920B94FDCEBEDBE803C0C849441220140A105C09163886";
    attribute INIT_35 of inst : label is "EFA7AFDF8EB4EF4D7F67557EE8EC7DB780E05440A023C0306E454944C26036BD";
    attribute INIT_36 of inst : label is "8F80FDC565940458E7FED9CB5E54FBAA9AE20B4234B428E90FBEC0D4F502C509";
    attribute INIT_37 of inst : label is "FDA7F51301B5BCEF7E83FF5B4A592EEF1BAAF2D8D39B684F1BA22A821107001A";
    attribute INIT_38 of inst : label is "3B0C820E201100248792E41252D92203F68FDFF87FBB63FFFFABF7D9ECCEBACD";
    attribute INIT_39 of inst : label is "3AA15608D3E08073A110421A41138838BF26493CB73F258EFA3CF96DFFA72FBE";
    attribute INIT_3A of inst : label is "61181930204008140A800389240C2220FBD73E37EF77A72D7DEDDD9EEBEFEFFB";
    attribute INIT_3B of inst : label is "148046C840A29B0EA2604E9D442EC026ACDC7FAB9FD2759CF7FEB1DDB7EFDE7F";
    attribute INIT_3C of inst : label is "DE9A083820034878414A218800371D057EE79F3FE8ED27FC9FBAEDF77A4F5F37";
    attribute INIT_3D of inst : label is "984118402578200F808308120026F7EE0EFA7BD69DE67E4D75FFBD8BEE75BEBF";
    attribute INIT_3E of inst : label is "2990C064A33A903598080002921904187FBEE1DC8BA5A7EFA4FE3EF35C6AFE6B";
    attribute INIT_3F of inst : label is "B0300C6004101029120690300B715011BEAEE97CFFADBF7DF796BF93D717FD7D";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "E19659E38E3871C38E19E591F9638E38E1D70EB87E4678EB8FFF400150580000";
    attribute INIT_01 of inst : label is "71C38E197E4659E38E38E1D70EB87F65919678EB8BAE1D70EB867919E3AE3870";
    attribute INIT_02 of inst : label is "679638E1C386591919E58E2E3871C38E19E4678E38E3875C3AE19E4678E38E38";
    attribute INIT_03 of inst : label is "9E4678EEBB875C3AE19E464678EB8B870E19679658E3870E19659678E3874E99";
    attribute INIT_04 of inst : label is "3875C3AE1FD9647E3AE2E3871C38E19E4678E38E1C38659659678EBB875C3AE1";
    attribute INIT_05 of inst : label is "8E2EB875C3AE19E4678E38E3871C38E19E47E38E38E1D70EB8659F1965F8E38E";
    attribute INIT_06 of inst : label is "1C38E19E4659E38E2E1C38679638E1D3A67D9638E9D3A659E58E3870E1967965";
    attribute INIT_07 of inst : label is "E1C386465919E58E38E1C70E38659F1919E38E38E1C70E387F6591FD8E38E387";
    attribute INIT_08 of inst : label is "59F1964638E1D3A679658E38E1D70EB87E464659678EB8E1C3865919679658E2";
    attribute INIT_09 of inst : label is "965F8E38C871C38E196597F65965F8E38E3875C3AE1F91FD918EB8B870E19646";
    attribute INIT_0A of inst : label is "9191F918E38E1D70EB87F659E3AE2E3871C38E19F647E38E38E1D70EB87F6591";
    attribute INIT_0B of inst : label is "E19F196597E38E2E3871C38E1967D919F638E38E1D70EB87F64659E38E3870E1";
    attribute INIT_0C of inst : label is "D965F8E38E3871C38E1965F919F658E38C871C38E1FD9191FC658E38E3871C38";
    attribute INIT_0D of inst : label is "E1D70EB87E596471FD8EE38E1D70EB867D965C764678EB8BAE1D70EB867965DD";
    attribute INIT_0E of inst : label is "E38E1C38659765DDD9E38B8E1C70E3867C7E38E38E1D70EB867C65919678EE38";
    attribute INIT_0F of inst : label is "8EAEB875C3AE19F765D91DD97E32B874E9FC6465D8E38E1C70E38659F647E5D8";
    attribute INIT_10 of inst : label is "2E1C386465919E58E3870E19196591F8E3870E197647E5D8E3874E997679771D";
    attribute INIT_11 of inst : label is "E19659678E3870E19191D971DDF8C870E1965979D965F8E3870E19665DFD918E";
    attribute INIT_12 of inst : label is "191964647E38E38E1C70E38679191DF8E38E3875C3AE1FDD91DDD91F8EB8B870";
    attribute INIT_13 of inst : label is "191FD97E4638E3870E19765D9F765DD8E2E1C3865D977E5D9638E3875C3AE1F9";
    attribute INIT_14 of inst : label is "EFBBFFC12FC17BC0000BAE1D70EB86791D9197E38EB874E997E4638E3871C38E";
    attribute INIT_15 of inst : label is "CCCDCDDCCCCCDCCDCCCDCDCCCDCCDCDCCDDDDDCDDDDCDDCCDCCCCCCCCCFABBEA";
    attribute INIT_16 of inst : label is "6B18D631AC652842528425084210865084B1AC6B1AD62FBEBBABFB9DDDCDDDCD";
    attribute INIT_17 of inst : label is "094A10C6B18C6B58CA52842504290852148CA52842108004010002065294A108";
    attribute INIT_18 of inst : label is "6B194A10942100080210040CA12942104214852908CA1284A18D631AC6318421";
    attribute INIT_19 of inst : label is "200840CA5084212942128421286528421294B58D6358D630842529421AC6B18C";
    attribute INIT_1A of inst : label is "358C631AC650842129410A5214852B29421284A0010042008194A10842120000";
    attribute INIT_1B of inst : label is "8431AC631AD6329421094A4200802008194A1084250C6358D6358CA5294A1096";
    attribute INIT_1C of inst : label is "8230A042815018D07110842A10AABFAAFEFACA50842129631AC631AC61084252";
    attribute INIT_1D of inst : label is "10A050350D468140A04429408506A10A0C6A140A506140A502810A88D28108C2";
    attribute INIT_1E of inst : label is "050210A84223408D2B41A20428140A5063450A04230A052234085062150846A1";
    attribute INIT_1F of inst : label is "518702C438CE118CE30E30906012C308CA18C251C210C25084A0B8A3F7F7D40A";
    attribute INIT_20 of inst : label is "1700C0300D4505540556880146388C7188E1C3218465186184238C671C230846";
    attribute INIT_21 of inst : label is "300E0581702C0B02E0180700C0300E0580601C0300E0180601C0300C03806018";
    attribute INIT_22 of inst : label is "241200882800AA0300C0302E0580601C0302E0580601C0B02C038060181700C0";
    attribute INIT_23 of inst : label is "000000000000000000AF54055154404051510140550000000004004558249248";
    attribute INIT_24 of inst : label is "0000000000000000042100000000000000000000000000001000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000002000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000010000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000800000000000000000000000000000040000000000000000000000";
    attribute INIT_28 of inst : label is "0000002000000000000004000000000000000000000000020000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000010842080000000000004000000000001000000";
    attribute INIT_2A of inst : label is "0008000000000000008008010040080004210820800000000000000000000000";
    attribute INIT_2B of inst : label is "4000800000400000000000100400820020000800000000800000000800020000";
    attribute INIT_2C of inst : label is "0108001004010040100401004010040100401004010802000400000010000000";
    attribute INIT_2D of inst : label is "0000000108200000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000401000200000000000040040001000000000000002000000000000000000";
    attribute INIT_2F of inst : label is "2108421000000842104100000000000000104000000104104200800100000000";
    attribute INIT_30 of inst : label is "4000000000000000000100000108400000000000000000000000000000001080";
    attribute INIT_31 of inst : label is "6FA24997274CED08400000000000000020000210800000000000000040000410";
    attribute INIT_32 of inst : label is "41EE286941BC2490A6420611111B845F4067B8DDEC90A485873C985D71C3BBBB";
    attribute INIT_33 of inst : label is "B9C713B52DBD96B39DC4BECF5F628FB6FB6FB67700035EE842850611111BB7C1";
    attribute INIT_34 of inst : label is "ABD7F7F7C4BFFFF2BDF59CE51DFAFCAA61A872B6D13235250690AE4FC049F624";
    attribute INIT_35 of inst : label is "59DDBD553E63DCA7AC64FCF27D72FE7A21C8498870308D13F0F274792CE299A5";
    attribute INIT_36 of inst : label is "F4C57F4D96DC7BB3EDBDE49C7F7F7F4F2811014A80AD1C00029592178053212B";
    attribute INIT_37 of inst : label is "9FBCF9FEABB1BF38F5E6CACF9FE0CF7D2C47353064E116A08418806454019826";
    attribute INIT_38 of inst : label is "FBE46A29282005A44900521DB8A8033BC76FBFABC07BFB9FABD4ADFA6C68D66D";
    attribute INIT_39 of inst : label is "4000110D977CB200054B261E09FE80B2FDAB2106FEF76D8B71C791E7FEE38DB3";
    attribute INIT_3A of inst : label is "0820328245442800D00004A4002E0340FFAE97FEF7FDFBFFF7CDFEFFFFD3F7B7";
    attribute INIT_3B of inst : label is "080400C02011006202E12A0520010048F6BF79FFBFBF7FF7AD7E1B3EF6FF7FD9";
    attribute INIT_3C of inst : label is "DD2E8C8F41278B08F485385CFAC585A0B4AD9E76B957EF1345F8BCEDE7BBDDBF";
    attribute INIT_3D of inst : label is "0AD044B101F845280008519B20866718D11CD87BDC3DC676D5F3BACB42D7ECB3";
    attribute INIT_3E of inst : label is "00340005000500095A303100001D000DE7FDFE7D9FAE7DFFDFFDFF7FFBC7FDBF";
    attribute INIT_3F of inst : label is "1046421082740400001110C210480041D4FE6EFDF7BAFBFFBF9FFF74FF4FEFDF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "408208A1041020810408A080A8210410408204102A0228410551501151100000";
    attribute INIT_01 of inst : label is "208104082A0208A10410408204102A20808228410904082041022808A1041020";
    attribute INIT_02 of inst : label is "228210408102080808A084241020810408A022841041020810408A0228410410";
    attribute INIT_03 of inst : label is "8A02284411020810408A02022841090204082282084102040820822841020408";
    attribute INIT_04 of inst : label is "102081040A88202A104241020810408A02284104081020820822841102081040";
    attribute INIT_05 of inst : label is "84241020810408A022841041020810408A02A1041040820410208A0820A84104";
    attribute INIT_06 of inst : label is "0810408A0208A10424081022821040810228821040810208A084102040822820";
    attribute INIT_07 of inst : label is "408102020808A0841040820410208A0808A10410408204102A2080A884104102";
    attribute INIT_08 of inst : label is "08A082021040810228208410408204102A020208228410408102080822820842";
    attribute INIT_09 of inst : label is "820A841040208104082082A20820A84104102081040A80A88084109020408202";
    attribute INIT_0A of inst : label is "8080A808410408204102A208A104241020810408A202A10410408204102A2080";
    attribute INIT_0B of inst : label is "408A082082A104241020810408228808A210410408204102A20208A104102040";
    attribute INIT_0C of inst : label is "8820A84104102081040820A808A208410402081040A88080A820841041020810";
    attribute INIT_0D of inst : label is "408204102A082020A88441040820410228820822022841090408204102282088";
    attribute INIT_0E of inst : label is "410408102082208888A1090408204102282A1041040820410228208082284410";
    attribute INIT_0F of inst : label is "84241020810408A2208808882A10102040A820208841040820410208A202A088";
    attribute INIT_10 of inst : label is "2408102020808A0841020408082080A8410204082202A0884102040822282208";
    attribute INIT_11 of inst : label is "40820822841020408080882088A84020408208288820A8410204082208A88084";
    attribute INIT_12 of inst : label is "080820202A10410408204102280808A84104102081040A888088880A84109020";
    attribute INIT_13 of inst : label is "080A882A02104102040822088A2208884240810208822A0882104102081040A8";
    attribute INIT_14 of inst : label is "40152AAA80002A800009040820410228088082A10410204082A0210410208104";
    attribute INIT_15 of inst : label is "5557467577656555554746547446565646746456576574765747464466405505";
    attribute INIT_16 of inst : label is "4A5294A5296108421084A5294A5296108425294A529490144115001676554674";
    attribute INIT_17 of inst : label is "0842101084210842C210842101084210842C2108421080842108421610842108";
    attribute INIT_18 of inst : label is "08584210842101084210842C210842101084210842C2108421294A5294A58421";
    attribute INIT_19 of inst : label is "294A52C210842108084210842161084210840421084210B08421084202108421";
    attribute INIT_1A of inst : label is "A5294A529610842108425294A5294B0842108421294A5294A5842108421094A5";
    attribute INIT_1B of inst : label is "8425294A5294B0842108421294A5294A5842108421094A5294A52C2108421084";
    attribute INIT_1C of inst : label is "8894A2528B454A513544A568944110140445C2108421084A5294A52961084210";
    attribute INIT_1D of inst : label is "44AA55344D568944AA556B44A552A94A2568955AD12B55A512894A2A528B5AD2";
    attribute INIT_1E of inst : label is "2D12B5A256A955A52B45A22528B44A5129445A252B5A252A945A512AB54AD289";
    attribute INIT_1F of inst : label is "538733C4784E308C611E1190E410C308CA184A11C650C6108CB5C57480A2144A";
    attribute INIT_20 of inst : label is "0B01401017EBBFAFEFA8A0005258847291E3C7109C2118E78C6384251C611842";
    attribute INIT_21 of inst : label is "503606813034050360280B0140D0160680A02C050160080202C050140580A008";
    attribute INIT_22 of inst : label is "241201555555FFFF0140D0360680A02C0D0360280A02C090040D80A0480B0340";
    attribute INIT_23 of inst : label is "000000000000000000EAFFBBAEBFAABEABFBFEAAFF000000000AAAEEF8249248";
    attribute INIT_24 of inst : label is "0000000000000000042100000000000000000000000000001000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000002000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000010000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000800000000000000000000000000000040000000000000000000000";
    attribute INIT_28 of inst : label is "0000002000000000000004000000000000000000000000020000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000010040080000000000004000000000001000000";
    attribute INIT_2A of inst : label is "0000000000000000000000010040080004010020000000000000000000000000";
    attribute INIT_2B of inst : label is "0010000000000000000000000000800000000000000000000000000000800000";
    attribute INIT_2C of inst : label is "0100000000000000000000000000000000000000010000000000000000000000";
    attribute INIT_2D of inst : label is "0000000108200000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000420000000000000000041000000000000000000002000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000004004000000000000000000000000000210000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000008020000000000000000000000000000001004";
    attribute INIT_31 of inst : label is "FD2012C403695108000000000000000000000010000000000000000000000010";
    attribute INIT_32 of inst : label is "95BB7E49894F0682B40A1E000003B0541402502A8E82B414B2C03AF64B95511F";
    attribute INIT_33 of inst : label is "D9EE775EFF94287A3A2B00208011600800800E090002094E02875E000003A9E0";
    attribute INIT_34 of inst : label is "53A5036B25C2FEC79AA1EC2E078CB53C2BFE91D297A7E19B26AAE597F47B69F9";
    attribute INIT_35 of inst : label is "97A63ABD1D65C2569BF774D4D88DC416B11BF3BEDD0F40484AA47EB9EB92A4E5";
    attribute INIT_36 of inst : label is "7BBD79FAF99DEFBF6EDBF3D6FEFFED3713121823EDA58189414AB3F26202F410";
    attribute INIT_37 of inst : label is "DB1DEF5FAD7FEFBEA3EC7BF5EBADABED0201698CC5D02970E2013803C002038D";
    attribute INIT_38 of inst : label is "C51E888DE504718C6E24688324201EBCC8DBF603CE3556BB7A7E5FA329B22766";
    attribute INIT_39 of inst : label is "41F522BEC8AC03423044AC5F48095B08D2C053F4F22F9747B773B62DD5D3A747";
    attribute INIT_3A of inst : label is "80A01380505002441C8AC008624080307FFBFFFFBEBBBDBF9F2EFEADEE6E7FAE";
    attribute INIT_3B of inst : label is "02200020821C1C044283C010A1410C61DB8EFFBFFFFAA3EFBDABFBAF9FFFFFEF";
    attribute INIT_3C of inst : label is "C304B1118E258A5741A08C48A3D4EE4A6DFB331DFB1DD9BC6FE9EDEB5BBEA5EF";
    attribute INIT_3D of inst : label is "000848144188122C5867002B127228E3C6FDFD377F9CD97CF34747FBABC2A747";
    attribute INIT_3E of inst : label is "045812A880C202013379012214084245FFBEFEA96FFB7FBFFFDE4F3EF6FFFEF9";
    attribute INIT_3F of inst : label is "80344400000040068840204451106043F53BD52DA3F56FFDCCFFFFEDFC5AF6E9";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000551450040400000";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000080000000000000000000000";
    attribute INIT_02 of inst : label is "0000000000000000000000200000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000080000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0000000000000000000200000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0020000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000200000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000000000000000000000002";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000000000000000008000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000200000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "0000000000000020000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000080000000000000000";
    attribute INIT_0E of inst : label is "0000000000000000000008000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0020000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "2000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000000000000008000";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000002000000000000000000000000000000";
    attribute INIT_14 of inst : label is "1101000000002A80000800000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "2023100221122022003301232123012300022022000320120022002000044554";
    attribute INIT_16 of inst : label is "5294A5294A4C6318C635294A5294A4C631A94A5294A501504541507220300003";
    attribute INIT_17 of inst : label is "6318C6210842108498C6318C6210842108498C6318C6310842108424C6318C63";
    attribute INIT_18 of inst : label is "109318C6318C6210842108498C6318C6210842108498C6318D4A5294A529318C";
    attribute INIT_19 of inst : label is "42108498C6318C6310842108424C6318C631884210842126318C6318C4210842";
    attribute INIT_1A of inst : label is "0842108424C6318C631884210842126318C6318C4210842109318C6318C62108";
    attribute INIT_1B of inst : label is "31884210842126318C6318C4210842109318C6318C6210842108498C6318C631";
    attribute INIT_1C of inst : label is "3319CC6711898CE27998C67138445105140498C6318C6310842108424C6318C6";
    attribute INIT_1D of inst : label is "98C4E2388E231188C4663198CE27119CCE31188C627188CE67319C4CE3338CE3";
    attribute INIT_1E of inst : label is "C66339C4E73388C67199CC4633198CE671988CCE338C4E33398C6673188C6711";
    attribute INIT_1F of inst : label is "1BCFA8E2BD6338C6B1AF3ACC751AE3BC671C6B78E378E758D6208A80A828998C";
    attribute INIT_20 of inst : label is "134350D42540511041460001035D56FAD577E3A9D6379C77C631C6B18EB18CE7";
    attribute INIT_21 of inst : label is "540680A1B4250D40684A134250142680A1A84D0141684A1A80D0941501A1A86A";
    attribute INIT_22 of inst : label is "008048000000AAAB4250140680A1A84D0140680A0A84D0141501A1280A034050";
    attribute INIT_23 of inst : label is "0000000000000000004004554015011150040000450000000005551101000001";
    attribute INIT_24 of inst : label is "0000000000000000040100000000000000000000000000001000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000002000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000010000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000800000000000000000000000000000040000000000000000000000";
    attribute INIT_28 of inst : label is "0000002000000000000004000000000000000000000000020000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000010040080000000000004000000000001000000";
    attribute INIT_2A of inst : label is "0000000000000000000000010040080004210820000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000800000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0100000000000000000000000000000000000000010000000000000000000000";
    attribute INIT_2D of inst : label is "0000000100200000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000400000000000000000040000000000000000000002000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000004100000000000000000000000000000200000000000000";
    attribute INIT_30 of inst : label is "4000000000000000000000000008400000000000000000000000000000001080";
    attribute INIT_31 of inst : label is "06C6DB436CADAE08400000000000000000000010800000000000000000000010";
    attribute INIT_32 of inst : label is "83826970810A8248912232BBBBBDA114A886127FF24892451044480A30AFFFF1";
    attribute INIT_33 of inst : label is "1C8A102A4DD2AB1703000000000000000000074C08888841888732BBBBBDA146";
    attribute INIT_34 of inst : label is "6F3FB3A819F56AB3ED77D985B6B1ACF9430F0E1442604428D47C4E21F210B800";
    attribute INIT_35 of inst : label is "FFEBE1E9F5F06F32D8F7A8DDBFBBBBED0495180770187218B2A044803242B354";
    attribute INIT_36 of inst : label is "87A5DFCEF3C4DD83003BDE2BED5E978EA1608A4E42430DC033A43589878763AB";
    attribute INIT_37 of inst : label is "8D035992E6594A48BF72AE1A05F2AFC5FC7305E6D0A0A1627E809C4E1BBFACCE";
    attribute INIT_38 of inst : label is "0068780209060018D480E0243E0020C9F9BF97FFDDFFD7FBF7525FB3F737DFFF";
    attribute INIT_39 of inst : label is "30000040820108D8BC19001045862906E59575BDD7BE7B4C56788DCDFDDDFFBF";
    attribute INIT_3A of inst : label is "9A93260146823469464488C201BBA25817B17F71DECEB85F9F9FFF7FEBDF3DF6";
    attribute INIT_3B of inst : label is "7371B924B60030A28411C0163950D4206DED6FEA9BF3DEBDB1CD3EF3EFFB875E";
    attribute INIT_3C of inst : label is "10E702480070002840843A90A2820416AFBFE75C5FD5BB3B5FFEA558BF79AFBD";
    attribute INIT_3D of inst : label is "10E70404056200820A031101021400475FE934FE79F77F6FE6E9BF77F4687FCD";
    attribute INIT_3E of inst : label is "04483891060A31183700618C960CA829EFFBE2F5F2F3DA476EFFD9EBD0633A7D";
    attribute INIT_3F of inst : label is "41520B9A89523CA0E49E715B000A01EAB612E33BFE3CBE1DDA335BD237FEF3FB";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000AABFBEBFFA00000";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000080000000000000000000000";
    attribute INIT_02 of inst : label is "0000000000000000000000200000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000080000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0000000000000000000200000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0020000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000200000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000000000000000000000002";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000000000000000008000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000200000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "0000000000000020000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000080000000000000000";
    attribute INIT_0E of inst : label is "0000000000000000000008000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0020000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "2000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000000000000008000";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000002000000000000000000000000000000";
    attribute INIT_14 of inst : label is "EEEAAAAAAAAA8000000800000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "02002300021103012300320102102301231103012310130123003312322EBFFB";
    attribute INIT_16 of inst : label is "084010840040000000000420080004001000210002002BEBFFAEBE8103032300";
    attribute INIT_17 of inst : label is "01084284A5084A1080000000284A5094A108000000001425284A508400008400";
    attribute INIT_18 of inst : label is "421000001084084A5094A1080020080084A10942108002108401080210810000";
    attribute INIT_19 of inst : label is "2942108000000000425084A508400000000021094A1084220004000012942129";
    attribute INIT_1A of inst : label is "252842508400000400021294A109420000020085094A129421000001004084A1";
    attribute INIT_1B of inst : label is "10A12942128420000000001084A508421000000084284A1094A1080000000014";
    attribute INIT_1C of inst : label is "A890AA42215448553000A42A90EEEEAFEAFE8000000000425084A50840000042";
    attribute INIT_1D of inst : label is "448855310C42A910885123548442A90AA4221548D52110AC42A9088056214842";
    attribute INIT_1E of inst : label is "A4429088520154846B10AAA4221548D521110AA42908856015484428910A4221";
    attribute INIT_1F of inst : label is "308710C438C6118C230E10886030C7184238C230C611C231843D5D55FFD5710A";
    attribute INIT_20 of inst : label is "0302409007FBABBFBBE8000002380C3180E1C3008461086184218C231C6118C2";
    attribute INIT_21 of inst : label is "9026068030140102606813034050260681200C050060681200C0D00401812048";
    attribute INIT_22 of inst : label is "000001555555FFFF014090060281204C050260280204C0D0240981A028130140";
    attribute INIT_23 of inst : label is "000000000000000000AEEFBFBFEAFEBEEFFBFFFFBA000000000AAAAAA0000000";
    attribute INIT_24 of inst : label is "0000000000000000040100000000000000000000000000001000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000002000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000010000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000800000000000000000000000000000040000000000000000000000";
    attribute INIT_28 of inst : label is "0000002000000000000004000000000000000000000000020000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000010040080000000000004000000000001000000";
    attribute INIT_2A of inst : label is "0000000000000000000000010040080004010020000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000800000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0100000000000000000000000000000000000000010000000000000000000000";
    attribute INIT_2D of inst : label is "0000000100200000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000400000000000000000040000000000000000000002000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000004000000000000000000000000000000200000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000008000000000000000000000000000000001000";
    attribute INIT_31 of inst : label is "884249C027C4CA08000000000000000000000010000000000000000000000010";
    attribute INIT_32 of inst : label is "A10A489101044600B00234333334A114AC4601555600B005D364506E012AAAA2";
    attribute INIT_33 of inst : label is "530F79FB6C9EB596EB000000000000000000061E0003880C888674333334A082";
    attribute INIT_34 of inst : label is "82E5D473C49817379FCBEDE5E75CEF2D1688A90197031388508104A0068A12A1";
    attribute INIT_35 of inst : label is "4B5F62DC61FB3CDB5FE7598FEADACB68136906D4A35E70190315881C41B832E1";
    attribute INIT_36 of inst : label is "8C423FFEDBF7CBDAAD68FCFFCDEBDA914F155A30663AE09218C5A41D26470837";
    attribute INIT_37 of inst : label is "E379F46B7E777344D9B507D1EA33FADA024E9452968A732D6608B840100E9050";
    attribute INIT_38 of inst : label is "A64200D2869210168711A68404227140CF7FFDF7FFFFA7BBD8FDBFBFFCACFFA7";
    attribute INIT_39 of inst : label is "AAE32B671E13CCC01078DA8699CD2086EF7577FD3F8BFFE2D7CA7F9FCCEFFFD7";
    attribute INIT_3A of inst : label is "4EAD662C94006284BD03C11404E608883BBF5DADFFFCCE27DE67FF9B4B96FDFB";
    attribute INIT_3B of inst : label is "2C8A29734C652880E22B2CE1C504FB082F0FD7EE79FBE7FFFAD6FA78F7F68EAA";
    attribute INIT_3C of inst : label is "63E42791C80E00809EC026C3232CC8516B8E41BF75D8BBFF7E55FCFBF37F9936";
    attribute INIT_3D of inst : label is "42A0490A1221243327472C803061AD68FE0FFFEBFEFB7FFFFEC7FEEDED8F6A34";
    attribute INIT_3E of inst : label is "91512405ACC3083180C3F00000047670BEB993CF1FD67FBFD4DAFABE5DBD79D7";
    attribute INIT_3F of inst : label is "AB048410220864C008C00DB6884D0081F42B59DF775FFAB6A51F2C2B751F5947";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
