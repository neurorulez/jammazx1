library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity splat_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of splat_sound is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CA",X"0F",X"8E",X"00",X"7F",X"CE",X"04",X"00",X"6F",X"01",X"6F",X"03",X"86",X"FF",X"A7",X"00",
		X"C6",X"80",X"E7",X"02",X"86",X"37",X"A7",X"03",X"86",X"3C",X"A7",X"01",X"E7",X"02",X"CE",X"00",
		X"7F",X"6F",X"00",X"09",X"26",X"FB",X"86",X"3C",X"97",X"01",X"0E",X"20",X"FE",X"7F",X"00",X"0B",
		X"97",X"09",X"36",X"CE",X"F1",X"49",X"A6",X"00",X"27",X"2D",X"7A",X"00",X"09",X"27",X"06",X"4C",
		X"BD",X"F1",X"1B",X"20",X"F1",X"08",X"DF",X"07",X"BD",X"F1",X"1B",X"DF",X"05",X"DE",X"07",X"A6",
		X"00",X"97",X"0E",X"A6",X"01",X"EE",X"02",X"DF",X"0C",X"8D",X"18",X"DE",X"07",X"08",X"08",X"08",
		X"08",X"DF",X"07",X"9C",X"05",X"26",X"E8",X"32",X"81",X"04",X"26",X"06",X"BD",X"F8",X"0D",X"7E",
		X"F8",X"73",X"39",X"CE",X"00",X"0F",X"81",X"00",X"27",X"15",X"81",X"03",X"27",X"09",X"C6",X"01",
		X"E7",X"00",X"08",X"80",X"02",X"20",X"EF",X"C6",X"91",X"E7",X"00",X"6F",X"01",X"08",X"08",X"C6",
		X"7E",X"E7",X"00",X"C6",X"F0",X"E7",X"01",X"C6",X"9D",X"E7",X"02",X"DE",X"0C",X"4F",X"F6",X"00",
		X"0A",X"5C",X"D7",X"0A",X"D4",X"0E",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",
		X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"54",X"89",X"00",X"48",X"48",X"48",X"48",X"48",
		X"B7",X"04",X"00",X"09",X"27",X"03",X"7E",X"00",X"0F",X"39",X"8E",X"00",X"7F",X"B6",X"04",X"02",
		X"43",X"8D",X"06",X"B6",X"04",X"02",X"0E",X"20",X"FE",X"84",X"1F",X"27",X"2D",X"81",X"06",X"2E",
		X"03",X"7E",X"F0",X"2D",X"0E",X"81",X"08",X"2E",X"05",X"80",X"07",X"7E",X"F7",X"C1",X"81",X"17",
		X"2E",X"08",X"80",X"09",X"BD",X"F8",X"0D",X"7E",X"F8",X"73",X"81",X"1F",X"2E",X"0C",X"80",X"18",
		X"CE",X"F1",X"0B",X"48",X"8D",X"15",X"EE",X"00",X"6E",X"00",X"39",X"FB",X"D7",X"FB",X"CC",X"FB",
		X"64",X"FB",X"C1",X"FB",X"EB",X"FC",X"10",X"F7",X"E7",X"FB",X"2F",X"DF",X"05",X"9B",X"06",X"97",
		X"06",X"96",X"05",X"89",X"00",X"97",X"05",X"DE",X"05",X"39",X"0F",X"8E",X"00",X"7F",X"CE",X"FF",
		X"FF",X"5F",X"E9",X"00",X"09",X"8C",X"F0",X"00",X"26",X"F8",X"E1",X"00",X"27",X"01",X"3E",X"86",
		X"04",X"BD",X"F8",X"0D",X"BD",X"F8",X"73",X"20",X"E1",X"30",X"6A",X"29",X"0A",X"AD",X"6A",X"0D",
		X"0E",X"41",X"00",X"29",X"01",X"55",X"6A",X"0D",X"0E",X"41",X"6A",X"29",X"0A",X"AD",X"00",X"29",
		X"01",X"55",X"6A",X"1D",X"05",X"FE",X"6A",X"29",X"05",X"56",X"6A",X"1D",X"05",X"FE",X"6A",X"0D",
		X"0E",X"41",X"6A",X"1D",X"05",X"FE",X"6A",X"29",X"05",X"56",X"3C",X"3C",X"04",X"0A",X"AA",X"00",
		X"04",X"02",X"AA",X"3C",X"04",X"0A",X"AA",X"00",X"04",X"02",X"AA",X"1E",X"3F",X"02",X"FE",X"3C",
		X"04",X"07",X"1C",X"3C",X"12",X"05",X"FA",X"3C",X"29",X"04",X"BE",X"3C",X"1D",X"05",X"53",X"3C",
		X"12",X"05",X"FA",X"00",X"12",X"02",X"3E",X"3C",X"12",X"05",X"FA",X"3C",X"1D",X"05",X"53",X"78",
		X"04",X"07",X"1C",X"3C",X"29",X"0E",X"3C",X"48",X"38",X"04",X"15",X"55",X"00",X"29",X"03",X"8F",
		X"38",X"04",X"0A",X"AA",X"1C",X"3F",X"05",X"FC",X"38",X"04",X"15",X"55",X"38",X"0D",X"09",X"80",
		X"38",X"12",X"08",X"F8",X"38",X"04",X"15",X"55",X"00",X"29",X"07",X"1E",X"38",X"04",X"0A",X"AA",
		X"00",X"0D",X"02",X"60",X"38",X"04",X"0A",X"AA",X"1C",X"1D",X"0F",X"FB",X"1C",X"29",X"07",X"1E",
		X"1C",X"30",X"06",X"B8",X"1C",X"3F",X"0B",X"F9",X"1C",X"30",X"06",X"B8",X"1C",X"29",X"07",X"1E",
		X"70",X"7C",X"04",X"05",X"55",X"00",X"0D",X"00",X"E4",X"7C",X"04",X"05",X"55",X"00",X"0D",X"00",
		X"E4",X"7C",X"04",X"05",X"55",X"00",X"04",X"01",X"FF",X"7C",X"1D",X"03",X"FE",X"00",X"12",X"00",
		X"D7",X"7C",X"12",X"04",X"7C",X"00",X"12",X"03",X"5D",X"7C",X"04",X"05",X"55",X"00",X"0D",X"00",
		X"E4",X"7C",X"04",X"05",X"55",X"00",X"0D",X"00",X"E4",X"7C",X"04",X"05",X"55",X"00",X"04",X"01",
		X"FF",X"7C",X"1D",X"03",X"FE",X"00",X"12",X"00",X"D7",X"7C",X"12",X"04",X"7C",X"00",X"12",X"03",
		X"5D",X"7C",X"04",X"05",X"55",X"00",X"0D",X"00",X"E4",X"7C",X"04",X"05",X"55",X"00",X"0D",X"00",
		X"E4",X"7C",X"04",X"05",X"55",X"7C",X"1D",X"03",X"FE",X"7C",X"12",X"04",X"7C",X"7C",X"29",X"05",
		X"56",X"98",X"F8",X"23",X"05",X"A8",X"F8",X"1D",X"05",X"FE",X"00",X"1D",X"02",X"FF",X"F8",X"17",
		X"06",X"59",X"F8",X"12",X"06",X"BA",X"00",X"12",X"0D",X"74",X"F8",X"0D",X"07",X"20",X"F8",X"09",
		X"07",X"8D",X"00",X"08",X"0F",X"1A",X"F8",X"0D",X"07",X"20",X"F8",X"17",X"06",X"59",X"00",X"0D",
		X"03",X"90",X"F8",X"0D",X"07",X"20",X"F8",X"08",X"07",X"8D",X"00",X"08",X"03",X"C6",X"7C",X"37",
		X"04",X"C1",X"7C",X"3F",X"04",X"7D",X"00",X"3F",X"02",X"3E",X"F8",X"1D",X"05",X"FE",X"F8",X"12",
		X"06",X"BA",X"00",X"12",X"03",X"5D",X"7C",X"37",X"04",X"C1",X"7C",X"3F",X"01",X"1F",X"7C",X"47",
		X"00",X"87",X"7C",X"3F",X"01",X"1F",X"7C",X"47",X"00",X"87",X"7C",X"3F",X"01",X"1F",X"7C",X"47",
		X"00",X"87",X"7C",X"3F",X"01",X"1F",X"7C",X"47",X"00",X"87",X"7C",X"3F",X"01",X"1F",X"7C",X"47",
		X"00",X"87",X"7C",X"3F",X"01",X"1F",X"7C",X"47",X"00",X"87",X"7C",X"3F",X"01",X"1F",X"7C",X"47",
		X"00",X"87",X"7C",X"3F",X"01",X"1F",X"7C",X"47",X"00",X"87",X"14",X"D4",X"1D",X"05",X"FE",X"D4",
		X"04",X"0F",X"FF",X"00",X"04",X"03",X"FF",X"6A",X"30",X"05",X"0A",X"D4",X"04",X"0F",X"FF",X"00",
		X"C6",X"03",X"D7",X"0B",X"4D",X"27",X"09",X"7C",X"00",X"0B",X"7C",X"00",X"0B",X"4A",X"20",X"F4",
		X"4F",X"B7",X"04",X"00",X"97",X"09",X"4F",X"91",X"09",X"26",X"03",X"73",X"04",X"00",X"D6",X"0B",
		X"5A",X"26",X"FD",X"4C",X"2A",X"F1",X"73",X"04",X"00",X"7C",X"00",X"09",X"2A",X"E8",X"39",X"C0",
		X"0D",X"37",X"BD",X"00",X"2C",X"33",X"C1",X"14",X"22",X"F5",X"01",X"96",X"24",X"9B",X"21",X"97",
		X"24",X"C9",X"F6",X"5A",X"2A",X"FD",X"96",X"28",X"4C",X"84",X"0F",X"8A",X"10",X"97",X"28",X"DE",
		X"27",X"E6",X"00",X"F7",X"04",X"00",X"84",X"0F",X"39",X"4F",X"CE",X"00",X"10",X"C6",X"61",X"A7",
		X"00",X"08",X"5A",X"26",X"FA",X"C6",X"5F",X"D7",X"26",X"C6",X"37",X"D7",X"30",X"C6",X"7E",X"D7",
		X"2C",X"CE",X"F5",X"64",X"DF",X"2D",X"D6",X"0C",X"D7",X"23",X"C0",X"03",X"BD",X"F3",X"56",X"08",
		X"D6",X"23",X"C0",X"02",X"BD",X"F3",X"4F",X"26",X"F7",X"D6",X"20",X"96",X"21",X"9B",X"0D",X"D9",
		X"0C",X"97",X"0D",X"D7",X"0C",X"DB",X"22",X"86",X"19",X"11",X"24",X"01",X"81",X"16",X"D7",X"23",
		X"01",X"C0",X"09",X"BD",X"F3",X"56",X"96",X"2F",X"16",X"48",X"C9",X"00",X"D7",X"2F",X"D6",X"23",
		X"C0",X"05",X"96",X"25",X"2A",X"06",X"7C",X"00",X"25",X"01",X"20",X"BE",X"5A",X"BD",X"F3",X"56",
		X"DE",X"0A",X"A6",X"00",X"2A",X"12",X"81",X"80",X"27",X"5F",X"4C",X"97",X"25",X"08",X"FF",X"00",
		X"0A",X"D6",X"23",X"C0",X"06",X"7E",X"F3",X"9A",X"08",X"E6",X"00",X"37",X"08",X"DF",X"0A",X"97",
		X"29",X"84",X"70",X"44",X"44",X"44",X"5F",X"8B",X"DD",X"C9",X"F4",X"97",X"2B",X"D7",X"2A",X"D6",
		X"23",X"D6",X"23",X"C0",X"0D",X"BD",X"F3",X"56",X"5F",X"DE",X"2A",X"EE",X"00",X"6E",X"00",X"96",
		X"29",X"47",X"C2",X"00",X"D4",X"0C",X"32",X"10",X"9B",X"0C",X"97",X"0C",X"08",X"D6",X"23",X"C0",
		X"0A",X"7E",X"F3",X"9C",X"96",X"29",X"47",X"C2",X"00",X"D4",X"22",X"32",X"10",X"9B",X"22",X"97",
		X"22",X"20",X"EA",X"32",X"DE",X"0A",X"09",X"6E",X"00",X"96",X"26",X"81",X"5F",X"2B",X"01",X"39",
		X"D6",X"23",X"C0",X"07",X"BD",X"F3",X"56",X"DE",X"25",X"6A",X"02",X"2B",X"12",X"EE",X"00",X"A6",
		X"00",X"36",X"08",X"DF",X"0A",X"F6",X"00",X"23",X"C0",X"09",X"BD",X"F3",X"56",X"20",X"55",X"EE",
		X"00",X"08",X"DF",X"0A",X"96",X"26",X"8B",X"03",X"97",X"26",X"D6",X"23",X"C0",X"07",X"01",X"7E",
		X"F3",X"9A",X"08",X"20",X"04",X"D7",X"20",X"D7",X"21",X"D6",X"29",X"C4",X"0F",X"CB",X"F8",X"C8",
		X"F8",X"32",X"9B",X"21",X"D9",X"20",X"97",X"21",X"D7",X"20",X"F6",X"00",X"23",X"C0",X"09",X"7E",
		X"F3",X"9A",X"96",X"26",X"80",X"03",X"97",X"26",X"DE",X"25",X"96",X"0B",X"D6",X"0A",X"8B",X"FF",
		X"C9",X"FF",X"E7",X"00",X"A7",X"01",X"D6",X"29",X"C4",X"0F",X"E7",X"02",X"D6",X"23",X"C0",X"0C",
		X"BD",X"F3",X"56",X"08",X"08",X"08",X"5F",X"01",X"32",X"47",X"49",X"C2",X"00",X"9B",X"0B",X"D9",
		X"0A",X"97",X"0B",X"F7",X"00",X"0A",X"D6",X"23",X"C0",X"07",X"7E",X"F3",X"9A",X"F4",X"1F",X"F4",
		X"34",X"F4",X"85",X"F4",X"82",X"F4",X"1F",X"F4",X"43",X"F4",X"A2",X"F4",X"C8",X"F6",X"61",X"F6",
		X"EA",X"F5",X"99",X"F6",X"92",X"F5",X"14",X"F6",X"A3",X"F5",X"3F",X"F5",X"D6",X"DE",X"2F",X"EE",
		X"03",X"08",X"DF",X"08",X"BD",X"F5",X"D0",X"08",X"39",X"EE",X"00",X"DF",X"08",X"CE",X"F5",X"D6",
		X"DF",X"2D",X"01",X"39",X"96",X"30",X"81",X"37",X"23",X"12",X"DE",X"2F",X"6A",X"02",X"2A",X"E9",
		X"80",X"03",X"97",X"30",X"CE",X"F4",X"FD",X"DF",X"2D",X"6D",X"00",X"39",X"CE",X"F5",X"34",X"DF",
		X"2D",X"01",X"20",X"05",X"08",X"08",X"01",X"8D",X"05",X"8D",X"03",X"6D",X"00",X"01",X"39",X"DE",
		X"2F",X"96",X"08",X"A7",X"03",X"96",X"09",X"A7",X"04",X"96",X"39",X"84",X"0F",X"A7",X"05",X"08",
		X"CE",X"F5",X"56",X"DF",X"2D",X"39",X"96",X"30",X"8B",X"03",X"97",X"30",X"CE",X"F5",X"D6",X"DF",
		X"2D",X"01",X"20",X"D5",X"7D",X"00",X"2F",X"26",X"CE",X"DE",X"08",X"A6",X"00",X"08",X"DF",X"08",
		X"97",X"39",X"2A",X"05",X"97",X"2F",X"A6",X"00",X"39",X"CE",X"F5",X"80",X"FF",X"00",X"2D",X"39",
		X"5F",X"96",X"39",X"84",X"70",X"44",X"44",X"44",X"8B",X"ED",X"C9",X"F4",X"D7",X"37",X"97",X"38",
		X"DE",X"37",X"EE",X"00",X"DF",X"2D",X"DF",X"2D",X"39",X"96",X"39",X"84",X"0F",X"4C",X"4C",X"97",
		X"2F",X"20",X"1D",X"7C",X"00",X"32",X"DE",X"31",X"8C",X"00",X"68",X"27",X"13",X"A6",X"00",X"CE",
		X"F5",X"EA",X"97",X"35",X"27",X"03",X"7E",X"F5",X"BC",X"CE",X"F5",X"A3",X"DF",X"2D",X"08",X"39",
		X"86",X"5E",X"B7",X"00",X"32",X"CE",X"F5",X"A3",X"7A",X"00",X"2F",X"27",X"03",X"7E",X"F5",X"D3",
		X"CE",X"F5",X"64",X"DF",X"2D",X"39",X"DE",X"08",X"5F",X"A6",X"00",X"4C",X"47",X"49",X"C2",X"00",
		X"9B",X"09",X"D9",X"08",X"97",X"09",X"D7",X"08",X"20",X"E6",X"96",X"32",X"80",X"5F",X"48",X"5F",
		X"9B",X"0F",X"D9",X"0E",X"D7",X"37",X"97",X"38",X"86",X"80",X"97",X"36",X"CE",X"F6",X"07",X"DF",
		X"2D",X"CE",X"00",X"10",X"DF",X"33",X"39",X"DE",X"37",X"EE",X"00",X"DF",X"37",X"CE",X"F6",X"1C",
		X"DF",X"2D",X"DE",X"31",X"A6",X"09",X"9B",X"35",X"A7",X"09",X"08",X"39",X"96",X"36",X"27",X"1D",
		X"74",X"00",X"36",X"DE",X"33",X"E6",X"00",X"94",X"37",X"26",X"09",X"FB",X"00",X"35",X"E7",X"00",
		X"7C",X"00",X"34",X"39",X"F0",X"00",X"35",X"E7",X"00",X"7C",X"00",X"34",X"39",X"D6",X"34",X"C1",
		X"20",X"27",X"0B",X"D6",X"38",X"D7",X"37",X"C6",X"80",X"F7",X"00",X"36",X"20",X"0F",X"CE",X"F5",
		X"64",X"D6",X"2F",X"26",X"03",X"7E",X"F6",X"5B",X"CE",X"F5",X"A3",X"DF",X"2D",X"6D",X"00",X"08",
		X"39",X"96",X"39",X"84",X"07",X"8B",X"60",X"97",X"32",X"DE",X"08",X"A6",X"00",X"08",X"DF",X"08",
		X"97",X"35",X"CE",X"F6",X"79",X"DF",X"2D",X"08",X"39",X"DE",X"31",X"5F",X"96",X"39",X"8B",X"F8",
		X"C2",X"00",X"E4",X"09",X"50",X"DB",X"35",X"D7",X"35",X"CE",X"F5",X"EA",X"DF",X"2D",X"08",X"08",
		X"01",X"39",X"D6",X"39",X"54",X"C4",X"07",X"CA",X"60",X"D7",X"32",X"C6",X"FF",X"C9",X"00",X"C9",
		X"00",X"20",X"E4",X"96",X"39",X"47",X"25",X"13",X"CE",X"00",X"00",X"DF",X"60",X"DF",X"62",X"DF",
		X"64",X"DF",X"66",X"08",X"CE",X"F5",X"64",X"FF",X"00",X"2D",X"39",X"85",X"02",X"26",X"0C",X"C6",
		X"5F",X"D7",X"32",X"CE",X"F6",X"D0",X"DF",X"2D",X"7E",X"F5",X"3B",X"FE",X"00",X"08",X"20",X"F6",
		X"5F",X"96",X"39",X"8B",X"AE",X"C2",X"00",X"D4",X"68",X"DE",X"08",X"A6",X"00",X"08",X"DF",X"08",
		X"10",X"97",X"35",X"CE",X"F5",X"EA",X"FF",X"00",X"2D",X"39",X"C6",X"60",X"D7",X"32",X"DE",X"08",
		X"E6",X"00",X"D7",X"37",X"08",X"DF",X"08",X"D6",X"39",X"54",X"24",X"18",X"CE",X"F7",X"2E",X"DF",
		X"2D",X"39",X"5F",X"96",X"38",X"47",X"C2",X"00",X"DE",X"31",X"E4",X"00",X"1B",X"A7",X"00",X"7C",
		X"00",X"32",X"A6",X"00",X"CE",X"F7",X"1A",X"DF",X"2D",X"39",X"78",X"00",X"37",X"25",X"13",X"27",
		X"06",X"7C",X"00",X"32",X"7E",X"F5",X"39",X"BD",X"F5",X"D0",X"6D",X"00",X"01",X"39",X"7A",X"00",
		X"32",X"08",X"A6",X"00",X"DE",X"08",X"A6",X"00",X"08",X"DF",X"08",X"97",X"38",X"CE",X"F7",X"02",
		X"DF",X"2D",X"39",X"00",X"00",X"55",X"55",X"33",X"33",X"25",X"DA",X"DA",X"25",X"C7",X"31",X"00",
		X"00",X"FF",X"FF",X"01",X"FE",X"53",X"00",X"66",X"16",X"66",X"1A",X"66",X"1E",X"66",X"21",X"66",
		X"24",X"08",X"FF",X"E2",X"66",X"1F",X"66",X"18",X"66",X"11",X"66",X"09",X"66",X"01",X"40",X"08",
		X"5A",X"08",X"00",X"FF",X"40",X"08",X"96",X"08",X"00",X"FF",X"40",X"08",X"C8",X"08",X"00",X"40",
		X"08",X"E6",X"08",X"00",X"40",X"08",X"FF",X"08",X"00",X"40",X"10",X"20",X"80",X"CC",X"CC",X"2F",
		X"80",X"E2",X"20",X"80",X"EC",X"2F",X"80",X"E2",X"20",X"80",X"EC",X"2F",X"80",X"E2",X"80",X"64",
		X"C4",X"80",X"53",X"00",X"08",X"05",X"0E",X"00",X"0D",X"05",X"FD",X"0D",X"00",X"0E",X"05",X"FD",
		X"70",X"F4",X"28",X"20",X"40",X"CE",X"20",X"00",X"80",X"F7",X"55",X"F7",X"8A",X"F7",X"A2",X"F7",
		X"B2",X"5F",X"D7",X"0D",X"48",X"48",X"8B",X"B9",X"C9",X"F7",X"D7",X"0A",X"97",X"0B",X"DE",X"0A",
		X"EE",X"00",X"DF",X"08",X"DE",X"0A",X"EE",X"02",X"E6",X"00",X"D7",X"0C",X"08",X"DF",X"0A",X"CE",
		X"F7",X"43",X"DF",X"0E",X"7E",X"F3",X"79",X"C6",X"BF",X"4F",X"B7",X"04",X"00",X"17",X"4A",X"26",
		X"FD",X"17",X"43",X"B7",X"04",X"00",X"8D",X"07",X"4A",X"26",X"FD",X"5A",X"26",X"EB",X"39",X"96",
		X"02",X"44",X"98",X"02",X"44",X"44",X"76",X"00",X"01",X"76",X"00",X"02",X"39",X"16",X"58",X"1B",
		X"1B",X"1B",X"CE",X"F9",X"F8",X"BD",X"F1",X"1B",X"A6",X"00",X"16",X"84",X"0F",X"97",X"0C",X"54",
		X"54",X"54",X"54",X"D7",X"0B",X"A6",X"01",X"16",X"54",X"54",X"54",X"54",X"D7",X"0D",X"84",X"0F",
		X"97",X"09",X"DF",X"03",X"CE",X"F9",X"40",X"7A",X"00",X"09",X"2B",X"08",X"A6",X"00",X"4C",X"BD",
		X"F1",X"1B",X"20",X"F3",X"DF",X"10",X"BD",X"F8",X"FF",X"DE",X"03",X"A6",X"02",X"97",X"12",X"BD",
		X"F9",X"11",X"DE",X"03",X"A6",X"03",X"97",X"0E",X"A6",X"04",X"97",X"0F",X"A6",X"05",X"16",X"A6",
		X"06",X"CE",X"FA",X"61",X"BD",X"F1",X"1B",X"17",X"DF",X"13",X"7F",X"00",X"1B",X"BD",X"F1",X"1B",
		X"DF",X"15",X"39",X"96",X"0B",X"97",X"1A",X"DE",X"13",X"DF",X"05",X"DE",X"05",X"A6",X"00",X"9B",
		X"1B",X"97",X"19",X"9C",X"15",X"27",X"26",X"D6",X"0C",X"08",X"DF",X"05",X"CE",X"00",X"1C",X"96",
		X"19",X"4A",X"26",X"FD",X"A6",X"00",X"B7",X"04",X"00",X"08",X"9C",X"17",X"26",X"F1",X"5A",X"27",
		X"DA",X"08",X"09",X"08",X"09",X"08",X"09",X"08",X"09",X"01",X"01",X"20",X"DF",X"96",X"0D",X"8D",
		X"60",X"7A",X"00",X"1A",X"26",X"C1",X"26",X"46",X"96",X"0E",X"27",X"42",X"7A",X"00",X"0F",X"27",
		X"3D",X"9B",X"1B",X"97",X"1B",X"DE",X"13",X"5F",X"96",X"1B",X"7D",X"00",X"0E",X"2B",X"06",X"AB",
		X"00",X"25",X"08",X"20",X"0B",X"AB",X"00",X"27",X"02",X"25",X"05",X"5D",X"27",X"08",X"20",X"0F",
		X"5D",X"26",X"03",X"DF",X"13",X"5C",X"08",X"9C",X"15",X"26",X"DD",X"5D",X"26",X"01",X"39",X"DF",
		X"15",X"96",X"0D",X"27",X"06",X"8D",X"08",X"96",X"12",X"8D",X"16",X"7E",X"F8",X"73",X"39",X"CE",
		X"00",X"1C",X"DF",X"07",X"DE",X"10",X"E6",X"00",X"08",X"BD",X"FB",X"1B",X"DE",X"07",X"DF",X"17",
		X"39",X"4D",X"27",X"2B",X"DE",X"10",X"DF",X"05",X"CE",X"00",X"1C",X"97",X"0A",X"DF",X"07",X"DE",
		X"05",X"D6",X"0A",X"D7",X"09",X"E6",X"01",X"54",X"54",X"54",X"54",X"08",X"DF",X"05",X"DE",X"07",
		X"A6",X"00",X"10",X"7A",X"00",X"09",X"26",X"FA",X"A7",X"00",X"08",X"9C",X"17",X"26",X"DE",X"39",
		X"08",X"7F",X"D9",X"FF",X"D9",X"7F",X"24",X"00",X"24",X"08",X"00",X"40",X"80",X"00",X"FF",X"00",
		X"80",X"40",X"10",X"7F",X"B0",X"D9",X"F5",X"FF",X"F5",X"D9",X"B0",X"7F",X"4E",X"24",X"09",X"00",
		X"09",X"24",X"4E",X"1C",X"80",X"40",X"29",X"1B",X"10",X"09",X"06",X"04",X"07",X"0C",X"12",X"1E",
		X"30",X"49",X"A4",X"C9",X"DF",X"EB",X"F6",X"FB",X"FF",X"FF",X"FB",X"F5",X"EA",X"DD",X"C7",X"9B",
		X"10",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",
		X"00",X"48",X"8A",X"95",X"A0",X"AB",X"B5",X"BF",X"C8",X"D1",X"DA",X"E1",X"E8",X"EE",X"F3",X"F7",
		X"FB",X"FD",X"FE",X"FF",X"FE",X"FD",X"FB",X"F7",X"F3",X"EE",X"E8",X"E1",X"DA",X"D1",X"C8",X"BF",
		X"B5",X"AB",X"A0",X"95",X"8A",X"7F",X"75",X"6A",X"5F",X"54",X"4A",X"40",X"37",X"2E",X"25",X"1E",
		X"17",X"11",X"0C",X"08",X"04",X"02",X"01",X"00",X"01",X"02",X"04",X"08",X"0C",X"11",X"17",X"1E",
		X"25",X"2E",X"37",X"40",X"4A",X"54",X"5F",X"6A",X"75",X"7F",X"0C",X"00",X"50",X"60",X"B0",X"20",
		X"20",X"F0",X"90",X"80",X"C0",X"50",X"70",X"10",X"7F",X"C5",X"EC",X"E7",X"BF",X"8D",X"6D",X"6A",
		X"7F",X"94",X"92",X"71",X"40",X"17",X"12",X"39",X"73",X"23",X"00",X"00",X"00",X"04",X"08",X"14",
		X"03",X"00",X"00",X"00",X"04",X"00",X"14",X"03",X"00",X"00",X"00",X"04",X"04",X"14",X"02",X"09",
		X"00",X"00",X"09",X"0C",X"11",X"02",X"00",X"00",X"00",X"28",X"15",X"1F",X"06",X"09",X"00",X"00",
		X"0F",X"3D",X"13",X"02",X"00",X"00",X"00",X"20",X"4C",X"11",X"02",X"00",X"00",X"00",X"18",X"15",
		X"15",X"02",X"05",X"00",X"00",X"16",X"6C",X"81",X"02",X"00",X"00",X"00",X"04",X"82",X"21",X"30",
		X"00",X"FF",X"00",X"1B",X"89",X"22",X"21",X"00",X"FE",X"00",X"1B",X"89",X"81",X"02",X"00",X"00",
		X"00",X"04",X"82",X"81",X"27",X"00",X"00",X"00",X"16",X"A4",X"68",X"20",X"00",X"02",X"26",X"03",
		X"86",X"20",X"18",X"20",X"01",X"01",X"30",X"28",X"30",X"08",X"10",X"20",X"30",X"20",X"10",X"0C",
		X"0A",X"08",X"07",X"06",X"05",X"04",X"60",X"45",X"28",X"21",X"5D",X"42",X"25",X"1E",X"58",X"3D",
		X"20",X"19",X"60",X"38",X"28",X"14",X"4C",X"31",X"14",X"0D",X"40",X"25",X"08",X"01",X"4C",X"31",
		X"14",X"0D",X"40",X"25",X"08",X"01",X"4C",X"31",X"14",X"0D",X"40",X"25",X"08",X"01",X"0A",X"09",
		X"08",X"07",X"06",X"05",X"06",X"07",X"08",X"09",X"0A",X"0A",X"0A",X"0A",X"0A",X"20",X"1F",X"1E",
		X"1D",X"1C",X"1B",X"1A",X"19",X"18",X"17",X"16",X"15",X"14",X"13",X"12",X"11",X"10",X"0F",X"0E",
		X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"07",X"06",X"05",X"05",X"05",X"05",X"05",X"1E",X"02",X"1B",
		X"04",X"23",X"07",X"1D",X"01",X"22",X"03",X"19",X"09",X"1F",X"06",X"1A",X"05",X"1C",X"0B",X"21",
		X"08",X"20",X"0A",X"60",X"45",X"28",X"21",X"03",X"04",X"24",X"01",X"01",X"02",X"02",X"04",X"04",
		X"08",X"08",X"10",X"10",X"30",X"60",X"C0",X"E0",X"01",X"01",X"02",X"02",X"03",X"04",X"05",X"06",
		X"07",X"08",X"09",X"0A",X"0C",X"01",X"01",X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"20",X"28",
		X"30",X"38",X"40",X"48",X"50",X"60",X"70",X"80",X"A0",X"B0",X"C0",X"36",X"A6",X"00",X"DF",X"05",
		X"DE",X"07",X"A7",X"00",X"08",X"DF",X"07",X"DE",X"05",X"08",X"5A",X"26",X"EF",X"32",X"39",X"86",
		X"01",X"97",X"13",X"C6",X"03",X"97",X"12",X"86",X"FF",X"B7",X"04",X"00",X"D7",X"0E",X"D6",X"0E",
		X"96",X"02",X"44",X"44",X"44",X"98",X"02",X"44",X"76",X"00",X"01",X"76",X"00",X"02",X"24",X"03",
		X"73",X"04",X"00",X"96",X"12",X"4A",X"26",X"FD",X"5A",X"26",X"E5",X"96",X"12",X"9B",X"13",X"97",
		X"12",X"26",X"DB",X"39",X"CE",X"FB",X"A3",X"DF",X"2D",X"DE",X"2D",X"A6",X"00",X"27",X"33",X"E6",
		X"01",X"C4",X"F0",X"D7",X"2C",X"E6",X"01",X"08",X"08",X"DF",X"2D",X"97",X"2B",X"C4",X"0F",X"96",
		X"2C",X"B7",X"04",X"00",X"96",X"2B",X"CE",X"00",X"05",X"09",X"26",X"FD",X"4A",X"26",X"F7",X"7F",
		X"04",X"00",X"96",X"2B",X"CE",X"00",X"05",X"09",X"26",X"FD",X"4A",X"26",X"F7",X"5A",X"26",X"DF",
		X"20",X"C7",X"39",X"01",X"FC",X"02",X"FC",X"03",X"F8",X"04",X"F8",X"06",X"F8",X"08",X"F4",X"0C",
		X"F4",X"10",X"F4",X"20",X"F2",X"40",X"F1",X"60",X"F1",X"80",X"F1",X"A0",X"F1",X"C0",X"F1",X"00",
		X"00",X"CE",X"FB",X"C7",X"7E",X"FC",X"5E",X"01",X"FF",X"01",X"00",X"10",X"CE",X"FB",X"D2",X"7E",
		X"FC",X"5E",X"80",X"F0",X"10",X"F0",X"06",X"CE",X"A5",X"00",X"DF",X"01",X"CE",X"FB",X"F1",X"BD",
		X"FD",X"40",X"CE",X"FC",X"01",X"BD",X"FC",X"49",X"7E",X"FC",X"E4",X"CE",X"FC",X"0B",X"7E",X"FC",
		X"5E",X"F0",X"10",X"03",X"20",X"34",X"B0",X"2A",X"02",X"18",X"40",X"70",X"30",X"02",X"0C",X"50",
		X"00",X"80",X"F0",X"20",X"01",X"01",X"18",X"F0",X"10",X"01",X"30",X"04",X"80",X"04",X"FE",X"30",
		X"CE",X"FC",X"06",X"8D",X"34",X"8D",X"14",X"8D",X"12",X"86",X"28",X"97",X"29",X"73",X"00",X"11",
		X"8D",X"3E",X"73",X"00",X"11",X"86",X"1E",X"8D",X"0D",X"20",X"EA",X"86",X"30",X"97",X"29",X"8D",
		X"2F",X"86",X"02",X"8D",X"01",X"39",X"16",X"CE",X"04",X"00",X"17",X"4A",X"26",X"FD",X"09",X"8C",
		X"00",X"00",X"26",X"F6",X"86",X"F0",X"97",X"0D",X"39",X"A6",X"00",X"97",X"24",X"A6",X"01",X"97",
		X"0D",X"A6",X"02",X"97",X"0C",X"A6",X"03",X"97",X"11",X"A6",X"04",X"97",X"29",X"39",X"8D",X"E9",
		X"8D",X"30",X"8D",X"58",X"96",X"28",X"91",X"29",X"26",X"F8",X"59",X"F7",X"04",X"00",X"8D",X"2D",
		X"8D",X"38",X"8D",X"5C",X"7D",X"00",X"0D",X"27",X"E4",X"7D",X"00",X"0E",X"26",X"E4",X"7D",X"00",
		X"11",X"27",X"DF",X"2B",X"05",X"7C",X"00",X"29",X"20",X"D8",X"7A",X"00",X"29",X"7A",X"00",X"28",
		X"20",X"D0",X"7F",X"00",X"0E",X"96",X"29",X"97",X"28",X"7F",X"00",X"27",X"39",X"96",X"02",X"44",
		X"44",X"44",X"98",X"02",X"97",X"22",X"08",X"84",X"07",X"39",X"96",X"22",X"44",X"76",X"00",X"01",
		X"76",X"00",X"02",X"86",X"00",X"24",X"02",X"96",X"0D",X"97",X"27",X"39",X"96",X"29",X"7A",X"00",
		X"28",X"27",X"04",X"08",X"09",X"20",X"08",X"97",X"28",X"D6",X"27",X"54",X"7C",X"00",X"0E",X"39",
		X"96",X"24",X"91",X"0E",X"27",X"04",X"08",X"09",X"20",X"09",X"7F",X"00",X"0E",X"96",X"0D",X"90",
		X"0C",X"97",X"0D",X"39",X"7F",X"00",X"1B",X"7F",X"00",X"25",X"86",X"0E",X"97",X"1C",X"7F",X"00",
		X"21",X"8D",X"9F",X"8D",X"A8",X"BD",X"FD",X"7A",X"8D",X"B0",X"BD",X"FD",X"7A",X"8D",X"BD",X"8D",
		X"79",X"8D",X"CD",X"8D",X"75",X"8D",X"0A",X"8D",X"71",X"8D",X"1D",X"8D",X"6D",X"8D",X"52",X"20",
		X"E2",X"96",X"20",X"7A",X"00",X"1C",X"27",X"07",X"B6",X"00",X"0D",X"26",X"0A",X"20",X"68",X"97",
		X"1C",X"96",X"1B",X"9B",X"25",X"97",X"1B",X"39",X"96",X"1B",X"91",X"23",X"27",X"07",X"08",X"96",
		X"0D",X"26",X"2A",X"20",X"29",X"7F",X"00",X"1B",X"7F",X"00",X"25",X"7F",X"00",X"21",X"DE",X"1D",
		X"A6",X"00",X"97",X"1A",X"27",X"17",X"A6",X"01",X"97",X"1F",X"A6",X"02",X"97",X"26",X"A6",X"03",
		X"97",X"20",X"A6",X"04",X"97",X"23",X"86",X"05",X"BD",X"F1",X"1B",X"DF",X"1D",X"39",X"32",X"32",
		X"39",X"96",X"1A",X"27",X"06",X"91",X"0D",X"26",X"04",X"20",X"03",X"08",X"09",X"39",X"7F",X"00",
		X"1A",X"96",X"1F",X"97",X"1B",X"96",X"26",X"97",X"25",X"39",X"96",X"21",X"9B",X"1B",X"97",X"21",
		X"2A",X"01",X"43",X"1B",X"B7",X"04",X"00",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"CA",X"F0",X"01",X"F1",X"2A",X"F0",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
