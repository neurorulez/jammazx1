library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity joust_sound is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of joust_sound is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"74",X"0F",X"8E",X"00",X"7F",X"CE",X"04",X"00",X"6F",X"01",X"6F",X"03",X"86",X"FF",X"A7",X"00",
		X"6F",X"02",X"86",X"37",X"A7",X"03",X"86",X"3C",X"A7",X"01",X"97",X"00",X"0E",X"20",X"FE",X"DF",
		X"07",X"CE",X"F0",X"C4",X"DF",X"02",X"86",X"80",X"D6",X"10",X"2A",X"09",X"D6",X"01",X"54",X"54",
		X"54",X"5C",X"5A",X"26",X"FD",X"7A",X"00",X"15",X"27",X"4C",X"7A",X"00",X"16",X"27",X"4C",X"7A",
		X"00",X"17",X"27",X"4C",X"7A",X"00",X"18",X"26",X"DF",X"D6",X"10",X"27",X"DB",X"C4",X"7F",X"D7",
		X"18",X"D6",X"01",X"58",X"DB",X"01",X"CB",X"0B",X"D7",X"01",X"7A",X"00",X"28",X"26",X"0E",X"D6",
		X"1C",X"D7",X"28",X"DE",X"02",X"09",X"8C",X"F0",X"BD",X"27",X"4E",X"DF",X"02",X"D6",X"01",X"2B",
		X"06",X"D4",X"14",X"C4",X"7F",X"20",X"05",X"D4",X"14",X"C4",X"7F",X"50",X"36",X"1B",X"16",X"32",
		X"DE",X"02",X"AD",X"00",X"20",X"A2",X"CE",X"00",X"0D",X"20",X"08",X"CE",X"00",X"0E",X"20",X"03",
		X"CE",X"00",X"0F",X"6D",X"18",X"27",X"12",X"6A",X"18",X"26",X"0E",X"E6",X"0C",X"E7",X"18",X"E6",
		X"00",X"EB",X"10",X"E1",X"14",X"27",X"12",X"E7",X"00",X"E6",X"00",X"E7",X"08",X"AB",X"04",X"60",
		X"04",X"16",X"DE",X"02",X"AD",X"00",X"7E",X"F0",X"28",X"DE",X"07",X"39",X"54",X"54",X"54",X"54",
		X"54",X"54",X"54",X"54",X"F7",X"04",X"00",X"39",X"CE",X"F2",X"9C",X"C6",X"1C",X"BD",X"F6",X"62",
		X"BD",X"F0",X"1F",X"39",X"CE",X"F2",X"F0",X"20",X"F2",X"CE",X"F3",X"0C",X"20",X"ED",X"86",X"80",
		X"97",X"10",X"86",X"F1",X"97",X"0E",X"86",X"80",X"97",X"0B",X"86",X"12",X"4A",X"26",X"FD",X"96",
		X"0D",X"9B",X"10",X"97",X"0D",X"44",X"44",X"44",X"8B",X"12",X"97",X"0F",X"DE",X"0E",X"A6",X"00",
		X"B7",X"04",X"00",X"7A",X"00",X"0B",X"26",X"E2",X"7A",X"00",X"10",X"96",X"10",X"81",X"20",X"26",
		X"D5",X"39",X"80",X"8C",X"98",X"A5",X"B0",X"BC",X"C6",X"D0",X"DA",X"E2",X"EA",X"F0",X"F5",X"FA",
		X"FD",X"FE",X"FF",X"FE",X"FD",X"FA",X"F5",X"F0",X"EA",X"E2",X"DA",X"D0",X"C6",X"BC",X"B0",X"A5",
		X"98",X"8C",X"80",X"73",X"67",X"5A",X"4F",X"43",X"39",X"2F",X"25",X"1D",X"15",X"0F",X"0A",X"05",
		X"02",X"01",X"00",X"01",X"02",X"05",X"0A",X"0F",X"15",X"1D",X"25",X"2F",X"39",X"43",X"4F",X"5A",
		X"67",X"73",X"7F",X"04",X"02",X"CE",X"F1",X"99",X"DF",X"0F",X"DE",X"0F",X"A6",X"00",X"27",X"33",
		X"E6",X"01",X"C4",X"F0",X"D7",X"0E",X"E6",X"01",X"08",X"08",X"DF",X"0F",X"97",X"0D",X"C4",X"0F",
		X"96",X"0E",X"B7",X"04",X"00",X"96",X"0D",X"CE",X"00",X"05",X"09",X"26",X"FD",X"4A",X"26",X"F7",
		X"7F",X"04",X"00",X"96",X"0D",X"CE",X"00",X"05",X"09",X"26",X"FD",X"4A",X"26",X"F7",X"5A",X"26",
		X"DF",X"20",X"C7",X"86",X"80",X"B7",X"04",X"02",X"39",X"01",X"FC",X"02",X"FC",X"03",X"F8",X"04",
		X"F8",X"06",X"F8",X"08",X"F4",X"0C",X"F4",X"10",X"F4",X"20",X"F2",X"40",X"F1",X"60",X"F1",X"80",
		X"F1",X"A0",X"F1",X"C0",X"F1",X"00",X"00",X"BD",X"F1",X"FA",X"BD",X"F2",X"13",X"39",X"CE",X"F3",
		X"82",X"20",X"F4",X"8D",X"F2",X"8D",X"27",X"20",X"FA",X"86",X"FF",X"97",X"04",X"CE",X"F3",X"9A",
		X"20",X"F1",X"C6",X"30",X"CE",X"F3",X"AC",X"8D",X"21",X"96",X"01",X"48",X"9B",X"01",X"8B",X"0B",
		X"97",X"01",X"44",X"44",X"8B",X"0C",X"97",X"0E",X"8D",X"29",X"5A",X"26",X"EC",X"39",X"96",X"04",
		X"80",X"08",X"2A",X"03",X"97",X"04",X"39",X"32",X"32",X"39",X"A6",X"00",X"97",X"0E",X"A6",X"01",
		X"97",X"0F",X"A6",X"02",X"97",X"10",X"A6",X"03",X"97",X"11",X"A6",X"04",X"97",X"12",X"A6",X"05",
		X"97",X"13",X"39",X"96",X"04",X"37",X"D6",X"12",X"D7",X"14",X"D6",X"0F",X"D7",X"15",X"43",X"D6",
		X"0E",X"B7",X"04",X"00",X"5A",X"26",X"FD",X"43",X"D6",X"0E",X"20",X"00",X"08",X"09",X"08",X"09",
		X"B7",X"04",X"00",X"5A",X"26",X"FD",X"7A",X"00",X"15",X"27",X"16",X"7A",X"00",X"14",X"26",X"DE",
		X"43",X"D6",X"12",X"B7",X"04",X"00",X"D7",X"14",X"D6",X"0E",X"9B",X"13",X"2B",X"1E",X"01",X"20",
		X"15",X"08",X"09",X"01",X"43",X"D6",X"0F",X"B7",X"04",X"00",X"D7",X"15",X"D6",X"0E",X"D0",X"10",
		X"D1",X"11",X"D1",X"11",X"27",X"06",X"D7",X"0E",X"C0",X"05",X"20",X"B8",X"33",X"39",X"DA",X"FF",
		X"DA",X"80",X"26",X"01",X"26",X"80",X"07",X"0A",X"07",X"00",X"F9",X"F6",X"F9",X"00",X"3A",X"3E",
		X"50",X"46",X"33",X"2C",X"27",X"20",X"25",X"1C",X"1A",X"17",X"14",X"11",X"10",X"33",X"08",X"03",
		X"02",X"01",X"02",X"03",X"04",X"05",X"06",X"0A",X"1E",X"32",X"70",X"00",X"FF",X"FF",X"FF",X"90",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"90",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"01",X"00",X"00",X"3F",X"3F",X"00",X"00",
		X"48",X"01",X"00",X"00",X"01",X"08",X"00",X"00",X"81",X"01",X"00",X"00",X"01",X"FF",X"00",X"00",
		X"01",X"08",X"00",X"00",X"01",X"10",X"00",X"00",X"3F",X"3F",X"00",X"00",X"01",X"10",X"00",X"00",
		X"05",X"05",X"00",X"00",X"01",X"01",X"00",X"00",X"31",X"FF",X"00",X"00",X"05",X"05",X"00",X"00",
		X"30",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"7F",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"04",X"00",X"00",X"04",
		X"7F",X"00",X"00",X"7F",X"04",X"00",X"00",X"04",X"FF",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"A0",X"0C",X"68",X"68",X"00",X"07",X"1F",X"0F",X"00",
		X"0C",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"01",X"04",X"00",X"00",X"3F",X"7F",X"00",X"00",X"01",X"04",X"00",X"00",
		X"05",X"FF",X"00",X"00",X"01",X"00",X"00",X"00",X"48",X"00",X"00",X"00",X"05",X"FF",X"00",X"00",
		X"02",X"80",X"00",X"30",X"0A",X"7F",X"00",X"7F",X"02",X"80",X"00",X"30",X"C0",X"80",X"00",X"20",
		X"01",X"10",X"00",X"15",X"C0",X"10",X"00",X"00",X"C0",X"80",X"00",X"00",X"FF",X"01",X"02",X"C3",
		X"FF",X"00",X"01",X"03",X"FF",X"80",X"FF",X"00",X"20",X"03",X"FF",X"50",X"FF",X"00",X"50",X"03",
		X"01",X"20",X"FF",X"00",X"FE",X"04",X"02",X"04",X"FF",X"00",X"48",X"03",X"01",X"0C",X"FF",X"00",
		X"48",X"02",X"01",X"0C",X"FF",X"00",X"E0",X"01",X"02",X"10",X"FF",X"00",X"50",X"FF",X"00",X"00",
		X"60",X"80",X"FF",X"02",X"01",X"06",X"FF",X"00",X"16",X"48",X"48",X"48",X"1B",X"CE",X"00",X"0D",
		X"DF",X"09",X"CE",X"F8",X"38",X"BD",X"F7",X"FA",X"C6",X"09",X"7E",X"F6",X"62",X"96",X"15",X"B7",
		X"04",X"00",X"96",X"0D",X"97",X"16",X"96",X"0E",X"97",X"17",X"DE",X"12",X"96",X"16",X"73",X"04",
		X"00",X"09",X"27",X"10",X"4A",X"26",X"FA",X"73",X"04",X"00",X"96",X"17",X"09",X"27",X"05",X"4A",
		X"26",X"FA",X"20",X"E8",X"B6",X"04",X"00",X"2B",X"01",X"43",X"8B",X"00",X"B7",X"04",X"00",X"96",
		X"16",X"9B",X"0F",X"97",X"16",X"96",X"17",X"9B",X"10",X"97",X"17",X"91",X"11",X"26",X"CB",X"96",
		X"14",X"27",X"06",X"9B",X"0D",X"97",X"0D",X"26",X"B9",X"39",X"CE",X"F4",X"20",X"7E",X"F4",X"CA",
		X"10",X"FF",X"01",X"01",X"01",X"CE",X"F4",X"44",X"DF",X"1E",X"BD",X"F5",X"AC",X"CE",X"A5",X"00",
		X"DF",X"00",X"CE",X"F4",X"6D",X"BD",X"F4",X"B5",X"BD",X"F5",X"50",X"CE",X"F4",X"72",X"BD",X"F4",
		X"B5",X"7E",X"F5",X"5D",X"90",X"10",X"02",X"14",X"40",X"B4",X"40",X"FF",X"14",X"30",X"D0",X"32",
		X"02",X"10",X"60",X"EE",X"20",X"02",X"08",X"54",X"E9",X"54",X"FF",X"20",X"28",X"C0",X"30",X"02",
		X"14",X"58",X"AC",X"20",X"02",X"08",X"58",X"A6",X"58",X"FF",X"18",X"22",X"00",X"30",X"10",X"FC",
		X"00",X"01",X"30",X"FC",X"01",X"00",X"01",X"10",X"F0",X"F0",X"01",X"30",X"CE",X"F4",X"77",X"8D",
		X"34",X"8D",X"14",X"8D",X"12",X"86",X"28",X"97",X"2A",X"73",X"00",X"12",X"8D",X"3E",X"73",X"00",
		X"12",X"86",X"1E",X"8D",X"0D",X"20",X"EA",X"86",X"30",X"97",X"2A",X"8D",X"2F",X"86",X"02",X"8D",
		X"01",X"39",X"16",X"CE",X"04",X"00",X"17",X"4A",X"26",X"FD",X"09",X"8C",X"00",X"00",X"26",X"F6",
		X"86",X"F0",X"97",X"0E",X"39",X"A6",X"00",X"97",X"25",X"A6",X"01",X"97",X"0E",X"A6",X"02",X"97",
		X"0D",X"A6",X"03",X"97",X"12",X"A6",X"04",X"97",X"2A",X"39",X"8D",X"E9",X"8D",X"30",X"8D",X"58",
		X"96",X"29",X"91",X"2A",X"26",X"F8",X"59",X"F7",X"04",X"00",X"8D",X"2D",X"8D",X"38",X"8D",X"5C",
		X"7D",X"00",X"0E",X"27",X"E4",X"7D",X"00",X"0F",X"26",X"E4",X"7D",X"00",X"12",X"27",X"DF",X"2B",
		X"05",X"7C",X"00",X"2A",X"20",X"D8",X"7A",X"00",X"2A",X"7A",X"00",X"29",X"20",X"D0",X"7F",X"00",
		X"0F",X"96",X"2A",X"97",X"29",X"7F",X"00",X"28",X"39",X"96",X"01",X"44",X"44",X"44",X"98",X"01",
		X"97",X"23",X"08",X"84",X"07",X"39",X"96",X"23",X"44",X"76",X"00",X"00",X"76",X"00",X"01",X"86",
		X"00",X"24",X"02",X"96",X"0E",X"97",X"28",X"39",X"96",X"2A",X"7A",X"00",X"29",X"27",X"04",X"08",
		X"09",X"20",X"08",X"97",X"29",X"D6",X"28",X"54",X"7C",X"00",X"0F",X"39",X"96",X"25",X"91",X"0F",
		X"27",X"04",X"08",X"09",X"20",X"09",X"7F",X"00",X"0F",X"96",X"0E",X"90",X"0D",X"97",X"0E",X"39",
		X"7F",X"00",X"1C",X"7F",X"00",X"26",X"86",X"0E",X"97",X"1D",X"7F",X"00",X"22",X"8D",X"9F",X"8D",
		X"A8",X"BD",X"F5",X"E6",X"8D",X"B0",X"BD",X"F5",X"E6",X"8D",X"BD",X"8D",X"79",X"8D",X"CD",X"8D",
		X"75",X"8D",X"0A",X"8D",X"71",X"8D",X"1D",X"8D",X"6D",X"8D",X"52",X"20",X"E2",X"96",X"21",X"7A",
		X"00",X"1D",X"27",X"07",X"B6",X"00",X"0E",X"26",X"0A",X"20",X"68",X"97",X"1D",X"96",X"1C",X"9B",
		X"26",X"97",X"1C",X"39",X"96",X"1C",X"91",X"24",X"27",X"07",X"08",X"96",X"0E",X"26",X"2A",X"20",
		X"29",X"7F",X"00",X"1C",X"7F",X"00",X"26",X"7F",X"00",X"22",X"DE",X"1E",X"A6",X"00",X"97",X"1B",
		X"27",X"17",X"A6",X"01",X"97",X"20",X"A6",X"02",X"97",X"27",X"A6",X"03",X"97",X"21",X"A6",X"04",
		X"97",X"24",X"86",X"05",X"BD",X"F7",X"FA",X"DF",X"1E",X"39",X"32",X"32",X"39",X"96",X"1B",X"27",
		X"06",X"91",X"0E",X"26",X"04",X"20",X"03",X"08",X"09",X"39",X"7F",X"00",X"1B",X"96",X"20",X"97",
		X"1C",X"96",X"27",X"97",X"26",X"39",X"96",X"22",X"9B",X"1C",X"97",X"22",X"2A",X"01",X"43",X"1B",
		X"B7",X"04",X"00",X"39",X"86",X"01",X"97",X"14",X"C6",X"03",X"20",X"00",X"97",X"13",X"86",X"FF",
		X"B7",X"04",X"00",X"D7",X"0F",X"D6",X"0F",X"96",X"01",X"44",X"44",X"44",X"98",X"01",X"44",X"76",
		X"00",X"00",X"76",X"00",X"01",X"24",X"03",X"73",X"04",X"00",X"96",X"13",X"4A",X"26",X"FD",X"5A",
		X"26",X"E5",X"96",X"13",X"9B",X"14",X"97",X"13",X"26",X"DB",X"39",X"97",X"0D",X"DF",X"10",X"D7",
		X"0E",X"D6",X"0F",X"96",X"01",X"44",X"44",X"44",X"98",X"01",X"44",X"76",X"00",X"00",X"76",X"00",
		X"01",X"86",X"00",X"24",X"02",X"96",X"0E",X"B7",X"04",X"00",X"DE",X"10",X"09",X"26",X"FD",X"5A",
		X"26",X"E1",X"D6",X"0E",X"D0",X"0D",X"27",X"09",X"DE",X"10",X"08",X"96",X"12",X"27",X"D0",X"20",
		X"CC",X"39",X"36",X"A6",X"00",X"DF",X"07",X"DE",X"09",X"A7",X"00",X"08",X"DF",X"09",X"DE",X"07",
		X"08",X"5A",X"26",X"EF",X"32",X"39",X"16",X"58",X"1B",X"1B",X"1B",X"CE",X"F9",X"27",X"BD",X"F7",
		X"FA",X"A6",X"00",X"16",X"84",X"0F",X"97",X"0E",X"54",X"54",X"54",X"54",X"D7",X"0D",X"A6",X"01",
		X"16",X"54",X"54",X"54",X"54",X"D7",X"0F",X"84",X"0F",X"97",X"0B",X"DF",X"05",X"CE",X"F8",X"38",
		X"7A",X"00",X"0B",X"2B",X"08",X"A6",X"00",X"4C",X"BD",X"F7",X"FA",X"20",X"F3",X"DF",X"12",X"BD",
		X"F7",X"68",X"DE",X"05",X"A6",X"02",X"97",X"14",X"BD",X"F7",X"7A",X"DE",X"05",X"A6",X"03",X"97",
		X"10",X"A6",X"04",X"97",X"11",X"A6",X"05",X"16",X"A6",X"06",X"CE",X"F9",X"BA",X"BD",X"F7",X"FA",
		X"17",X"DF",X"15",X"7F",X"00",X"1D",X"BD",X"F7",X"FA",X"DF",X"17",X"39",X"96",X"0D",X"97",X"1C",
		X"DE",X"15",X"DF",X"07",X"DE",X"07",X"A6",X"00",X"9B",X"1D",X"97",X"1B",X"9C",X"17",X"27",X"26",
		X"D6",X"0E",X"08",X"DF",X"07",X"CE",X"00",X"1E",X"96",X"1B",X"4A",X"26",X"FD",X"A6",X"00",X"B7",
		X"04",X"00",X"08",X"9C",X"19",X"26",X"F1",X"5A",X"27",X"DA",X"08",X"09",X"08",X"09",X"08",X"09",
		X"08",X"09",X"01",X"01",X"20",X"DF",X"96",X"0F",X"8D",X"60",X"7A",X"00",X"1C",X"26",X"C1",X"26",
		X"46",X"96",X"10",X"27",X"42",X"7A",X"00",X"11",X"27",X"3D",X"9B",X"1D",X"97",X"1D",X"DE",X"15",
		X"5F",X"96",X"1D",X"7D",X"00",X"10",X"2B",X"06",X"AB",X"00",X"25",X"08",X"20",X"0B",X"AB",X"00",
		X"27",X"02",X"25",X"05",X"5D",X"27",X"08",X"20",X"0F",X"5D",X"26",X"03",X"DF",X"15",X"5C",X"08",
		X"9C",X"17",X"26",X"DD",X"5D",X"26",X"01",X"39",X"DF",X"17",X"96",X"0F",X"27",X"06",X"8D",X"08",
		X"96",X"14",X"8D",X"16",X"7E",X"F6",X"DC",X"39",X"CE",X"00",X"1E",X"DF",X"09",X"DE",X"12",X"E6",
		X"00",X"08",X"BD",X"F6",X"62",X"DE",X"09",X"DF",X"19",X"39",X"4D",X"27",X"2B",X"DE",X"12",X"DF",
		X"07",X"CE",X"00",X"1E",X"97",X"0C",X"DF",X"09",X"DE",X"07",X"D6",X"0C",X"D7",X"0B",X"E6",X"01",
		X"54",X"54",X"54",X"54",X"08",X"DF",X"07",X"DE",X"09",X"A6",X"00",X"10",X"7A",X"00",X"0B",X"26",
		X"FA",X"A7",X"00",X"08",X"9C",X"19",X"26",X"DE",X"39",X"8E",X"00",X"7F",X"B6",X"04",X"02",X"CE",
		X"F0",X"C4",X"DF",X"02",X"CE",X"00",X"0D",X"DF",X"09",X"C6",X"AF",X"D7",X"04",X"0E",X"43",X"84",
		X"3F",X"4D",X"27",X"34",X"4A",X"81",X"14",X"22",X"08",X"BD",X"F6",X"76",X"BD",X"F6",X"DC",X"20",
		X"27",X"81",X"1F",X"22",X"0F",X"80",X"15",X"CE",X"F8",X"22",X"48",X"BD",X"F7",X"FA",X"EE",X"00",
		X"AD",X"00",X"20",X"14",X"81",X"22",X"22",X"07",X"80",X"20",X"BD",X"FF",X"4A",X"20",X"09",X"81",
		X"26",X"22",X"05",X"80",X"23",X"BD",X"FF",X"6C",X"20",X"FE",X"DF",X"07",X"9B",X"08",X"97",X"08",
		X"24",X"03",X"7C",X"00",X"07",X"DE",X"07",X"39",X"0F",X"8E",X"00",X"7F",X"CE",X"FF",X"FF",X"5F",
		X"E9",X"00",X"09",X"8C",X"F0",X"00",X"26",X"F8",X"E1",X"00",X"27",X"01",X"3E",X"BD",X"F1",X"52",
		X"20",X"E6",X"F5",X"F4",X"F0",X"D4",X"F0",X"D9",X"F0",X"C8",X"F1",X"BE",X"F1",X"C9",X"F1",X"D2",
		X"F1",X"52",X"F0",X"DE",X"F0",X"01",X"FF",X"44",X"08",X"7F",X"D9",X"FF",X"D9",X"7F",X"24",X"00",
		X"24",X"08",X"00",X"40",X"80",X"00",X"FF",X"00",X"80",X"40",X"10",X"7F",X"B0",X"D9",X"F5",X"FF",
		X"F5",X"D9",X"B0",X"7F",X"4E",X"24",X"09",X"00",X"09",X"24",X"4E",X"10",X"7F",X"C5",X"EC",X"E7",
		X"BF",X"8D",X"6D",X"6A",X"7F",X"94",X"92",X"71",X"40",X"17",X"12",X"39",X"10",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"48",X"8A",X"95",
		X"A0",X"AB",X"B5",X"BF",X"C8",X"D1",X"DA",X"E1",X"E8",X"EE",X"F3",X"F7",X"FB",X"FD",X"FE",X"FF",
		X"FE",X"FD",X"FB",X"F7",X"F3",X"EE",X"E8",X"E1",X"DA",X"D1",X"C8",X"BF",X"B5",X"AB",X"A0",X"95",
		X"8A",X"7F",X"75",X"6A",X"5F",X"54",X"4A",X"40",X"37",X"2E",X"25",X"1E",X"17",X"11",X"0C",X"08",
		X"04",X"02",X"01",X"00",X"01",X"02",X"04",X"08",X"0C",X"11",X"17",X"1E",X"25",X"2E",X"37",X"40",
		X"4A",X"54",X"5F",X"6A",X"75",X"7F",X"10",X"59",X"7B",X"98",X"AC",X"B3",X"AC",X"98",X"7B",X"59",
		X"37",X"19",X"06",X"00",X"06",X"19",X"37",X"08",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"10",X"76",X"FF",X"B8",X"D0",X"9D",X"E6",X"6A",X"82",X"76",X"EA",X"81",X"86",X"4E",X"9C",X"32",
		X"63",X"10",X"00",X"F4",X"00",X"E8",X"00",X"DC",X"00",X"E2",X"00",X"DC",X"00",X"E8",X"00",X"F4",
		X"00",X"00",X"24",X"7F",X"B0",X"D6",X"E8",X"E3",X"C9",X"A3",X"7B",X"5E",X"54",X"5E",X"7B",X"A3",
		X"C9",X"E3",X"E8",X"D6",X"B0",X"7F",X"4C",X"26",X"14",X"19",X"33",X"5A",X"81",X"9E",X"A8",X"9E",
		X"81",X"5A",X"33",X"19",X"14",X"26",X"4C",X"11",X"05",X"11",X"01",X"0F",X"01",X"3A",X"21",X"35",
		X"11",X"FF",X"00",X"0D",X"0E",X"15",X"00",X"00",X"FD",X"00",X"01",X"4E",X"31",X"11",X"00",X"01",
		X"00",X"03",X"4F",X"F6",X"53",X"03",X"00",X"02",X"06",X"79",X"14",X"17",X"00",X"00",X"00",X"0E",
		X"00",X"13",X"10",X"00",X"FF",X"00",X"09",X"80",X"F2",X"19",X"00",X"00",X"00",X"16",X"8F",X"41",
		X"02",X"D0",X"00",X"00",X"27",X"52",X"52",X"36",X"00",X"00",X"00",X"10",X"24",X"73",X"29",X"03",
		X"00",X"00",X"10",X"A6",X"11",X"40",X"03",X"ED",X"09",X"09",X"1B",X"16",X"82",X"03",X"0E",X"01",
		X"0E",X"7F",X"11",X"29",X"00",X"F0",X"05",X"08",X"B6",X"63",X"26",X"06",X"00",X"00",X"10",X"A6",
		X"21",X"25",X"00",X"03",X"0A",X"03",X"4F",X"43",X"0A",X"00",X"04",X"02",X"0D",X"0E",X"1F",X"12",
		X"00",X"FF",X"10",X"04",X"4E",X"11",X"10",X"00",X"0A",X"00",X"01",X"80",X"21",X"30",X"00",X"FF",
		X"00",X"1B",X"00",X"22",X"21",X"00",X"FE",X"00",X"1B",X"00",X"01",X"01",X"02",X"02",X"04",X"04",
		X"08",X"08",X"10",X"10",X"30",X"60",X"C0",X"E0",X"01",X"01",X"02",X"02",X"03",X"04",X"05",X"06",
		X"07",X"08",X"09",X"0A",X"0C",X"80",X"7C",X"78",X"74",X"70",X"74",X"78",X"7C",X"80",X"01",X"01",
		X"02",X"02",X"04",X"04",X"08",X"08",X"10",X"20",X"28",X"30",X"38",X"40",X"48",X"50",X"60",X"70",
		X"80",X"A0",X"B0",X"C0",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",
		X"08",X"40",X"08",X"40",X"08",X"40",X"08",X"40",X"40",X"10",X"08",X"01",X"01",X"01",X"01",X"01",
		X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"06",X"08",X"0A",X"0C",X"10",X"14",X"18",X"20",X"30",
		X"40",X"50",X"40",X"30",X"20",X"10",X"0C",X"0A",X"08",X"07",X"06",X"05",X"04",X"03",X"02",X"02",
		X"01",X"01",X"01",X"07",X"08",X"09",X"0A",X"0C",X"08",X"0C",X"08",X"80",X"10",X"78",X"18",X"70",
		X"20",X"60",X"28",X"58",X"30",X"50",X"40",X"48",X"00",X"01",X"40",X"02",X"42",X"03",X"43",X"04",
		X"44",X"05",X"45",X"06",X"46",X"07",X"47",X"08",X"48",X"09",X"49",X"0A",X"4A",X"0B",X"4B",X"00",
		X"14",X"18",X"20",X"30",X"40",X"50",X"40",X"30",X"20",X"10",X"0C",X"0A",X"08",X"07",X"06",X"05",
		X"CC",X"BB",X"60",X"10",X"EE",X"AA",X"50",X"00",X"28",X"43",X"29",X"31",X"39",X"38",X"32",X"20",
		X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",
		X"4E",X"49",X"43",X"53",X"C0",X"0D",X"37",X"BD",X"00",X"2C",X"33",X"C1",X"14",X"22",X"F5",X"01",
		X"96",X"24",X"9B",X"21",X"97",X"24",X"C9",X"F6",X"5A",X"2A",X"FD",X"96",X"28",X"4C",X"84",X"0F",
		X"8A",X"10",X"97",X"28",X"DE",X"27",X"E6",X"00",X"F7",X"04",X"00",X"84",X"0F",X"39",X"4F",X"CE",
		X"00",X"10",X"C6",X"61",X"A7",X"00",X"08",X"5A",X"26",X"FA",X"C6",X"5F",X"D7",X"26",X"C6",X"37",
		X"D7",X"30",X"C6",X"7E",X"D7",X"2C",X"CE",X"FC",X"A9",X"DF",X"2D",X"D6",X"0C",X"D7",X"23",X"C0",
		X"03",X"BD",X"FA",X"9B",X"08",X"D6",X"23",X"C0",X"02",X"BD",X"FA",X"94",X"26",X"F7",X"D6",X"20",
		X"96",X"21",X"9B",X"0D",X"D9",X"0C",X"97",X"0D",X"D7",X"0C",X"DB",X"22",X"86",X"19",X"11",X"24",
		X"01",X"81",X"16",X"D7",X"23",X"01",X"C0",X"09",X"BD",X"FA",X"9B",X"96",X"2F",X"16",X"48",X"C9",
		X"00",X"D7",X"2F",X"D6",X"23",X"C0",X"05",X"96",X"25",X"2A",X"06",X"7C",X"00",X"25",X"01",X"20",
		X"BE",X"5A",X"BD",X"FA",X"9B",X"DE",X"0A",X"A6",X"00",X"2A",X"12",X"81",X"80",X"27",X"5F",X"4C",
		X"97",X"25",X"08",X"FF",X"00",X"0A",X"D6",X"23",X"C0",X"06",X"7E",X"FA",X"DF",X"08",X"E6",X"00",
		X"37",X"08",X"DF",X"0A",X"97",X"29",X"84",X"70",X"44",X"44",X"44",X"5F",X"8B",X"22",X"C9",X"FC",
		X"97",X"2B",X"D7",X"2A",X"D6",X"23",X"D6",X"23",X"C0",X"0D",X"BD",X"FA",X"9B",X"5F",X"DE",X"2A",
		X"EE",X"00",X"6E",X"00",X"96",X"29",X"47",X"C2",X"00",X"D4",X"0C",X"32",X"10",X"9B",X"0C",X"97",
		X"0C",X"08",X"D6",X"23",X"C0",X"0A",X"7E",X"FA",X"E1",X"96",X"29",X"47",X"C2",X"00",X"D4",X"22",
		X"32",X"10",X"9B",X"22",X"97",X"22",X"20",X"EA",X"32",X"DE",X"0A",X"09",X"6E",X"00",X"96",X"26",
		X"81",X"5F",X"2B",X"01",X"39",X"D6",X"23",X"C0",X"07",X"BD",X"FA",X"9B",X"DE",X"25",X"6A",X"02",
		X"2B",X"12",X"EE",X"00",X"A6",X"00",X"36",X"08",X"DF",X"0A",X"F6",X"00",X"23",X"C0",X"09",X"BD",
		X"FA",X"9B",X"20",X"55",X"EE",X"00",X"08",X"DF",X"0A",X"96",X"26",X"8B",X"03",X"97",X"26",X"D6",
		X"23",X"C0",X"07",X"01",X"7E",X"FA",X"DF",X"08",X"20",X"04",X"D7",X"20",X"D7",X"21",X"D6",X"29",
		X"C4",X"0F",X"CB",X"F8",X"C8",X"F8",X"32",X"9B",X"21",X"D9",X"20",X"97",X"21",X"D7",X"20",X"F6",
		X"00",X"23",X"C0",X"09",X"7E",X"FA",X"DF",X"96",X"26",X"80",X"03",X"97",X"26",X"DE",X"25",X"96",
		X"0B",X"D6",X"0A",X"8B",X"FF",X"C9",X"FF",X"E7",X"00",X"A7",X"01",X"D6",X"29",X"C4",X"0F",X"E7",
		X"02",X"D6",X"23",X"C0",X"0C",X"BD",X"FA",X"9B",X"08",X"08",X"08",X"5F",X"01",X"32",X"47",X"49",
		X"C2",X"00",X"9B",X"0B",X"D9",X"0A",X"97",X"0B",X"F7",X"00",X"0A",X"D6",X"23",X"C0",X"07",X"7E",
		X"FA",X"DF",X"FB",X"64",X"FB",X"79",X"FB",X"CA",X"FB",X"C7",X"FB",X"64",X"FB",X"88",X"FB",X"E7",
		X"FC",X"0D",X"FD",X"A6",X"FE",X"2F",X"FC",X"DE",X"FD",X"D7",X"FC",X"59",X"FD",X"E8",X"FC",X"84",
		X"FD",X"1B",X"DE",X"2F",X"EE",X"03",X"08",X"DF",X"08",X"BD",X"FD",X"15",X"08",X"39",X"EE",X"00",
		X"DF",X"08",X"CE",X"FD",X"1B",X"DF",X"2D",X"01",X"39",X"96",X"30",X"81",X"37",X"23",X"12",X"DE",
		X"2F",X"6A",X"02",X"2A",X"E9",X"80",X"03",X"97",X"30",X"CE",X"FC",X"42",X"DF",X"2D",X"6D",X"00",
		X"39",X"CE",X"FC",X"79",X"DF",X"2D",X"01",X"20",X"05",X"08",X"08",X"01",X"8D",X"05",X"8D",X"03",
		X"6D",X"00",X"01",X"39",X"DE",X"2F",X"96",X"08",X"A7",X"03",X"96",X"09",X"A7",X"04",X"96",X"39",
		X"84",X"0F",X"A7",X"05",X"08",X"CE",X"FC",X"9B",X"DF",X"2D",X"39",X"96",X"30",X"8B",X"03",X"97",
		X"30",X"CE",X"FD",X"1B",X"DF",X"2D",X"01",X"20",X"D5",X"7D",X"00",X"2F",X"26",X"CE",X"DE",X"08",
		X"A6",X"00",X"08",X"DF",X"08",X"97",X"39",X"2A",X"05",X"97",X"2F",X"A6",X"00",X"39",X"CE",X"FC",
		X"C5",X"FF",X"00",X"2D",X"39",X"5F",X"96",X"39",X"84",X"70",X"44",X"44",X"44",X"8B",X"32",X"C9",
		X"FC",X"D7",X"37",X"97",X"38",X"DE",X"37",X"EE",X"00",X"DF",X"2D",X"DF",X"2D",X"39",X"96",X"39",
		X"84",X"0F",X"4C",X"4C",X"97",X"2F",X"20",X"1D",X"7C",X"00",X"32",X"DE",X"31",X"8C",X"00",X"68",
		X"27",X"13",X"A6",X"00",X"CE",X"FD",X"2F",X"97",X"35",X"27",X"03",X"7E",X"FD",X"01",X"CE",X"FC",
		X"E8",X"DF",X"2D",X"08",X"39",X"86",X"5E",X"B7",X"00",X"32",X"CE",X"FC",X"E8",X"7A",X"00",X"2F",
		X"27",X"03",X"7E",X"FD",X"18",X"CE",X"FC",X"A9",X"DF",X"2D",X"39",X"DE",X"08",X"5F",X"A6",X"00",
		X"4C",X"47",X"49",X"C2",X"00",X"9B",X"09",X"D9",X"08",X"97",X"09",X"D7",X"08",X"20",X"E6",X"96",
		X"32",X"80",X"5F",X"48",X"5F",X"9B",X"0F",X"D9",X"0E",X"D7",X"37",X"97",X"38",X"86",X"80",X"97",
		X"36",X"CE",X"FD",X"4C",X"DF",X"2D",X"CE",X"00",X"10",X"DF",X"33",X"39",X"DE",X"37",X"EE",X"00",
		X"DF",X"37",X"CE",X"FD",X"61",X"DF",X"2D",X"DE",X"31",X"A6",X"09",X"9B",X"35",X"A7",X"09",X"08",
		X"39",X"96",X"36",X"27",X"1D",X"74",X"00",X"36",X"DE",X"33",X"E6",X"00",X"94",X"37",X"26",X"09",
		X"FB",X"00",X"35",X"E7",X"00",X"7C",X"00",X"34",X"39",X"F0",X"00",X"35",X"E7",X"00",X"7C",X"00",
		X"34",X"39",X"D6",X"34",X"C1",X"20",X"27",X"0B",X"D6",X"38",X"D7",X"37",X"C6",X"80",X"F7",X"00",
		X"36",X"20",X"0F",X"CE",X"FC",X"A9",X"D6",X"2F",X"26",X"03",X"7E",X"FD",X"A0",X"CE",X"FC",X"E8",
		X"DF",X"2D",X"6D",X"00",X"08",X"39",X"96",X"39",X"84",X"07",X"8B",X"60",X"97",X"32",X"DE",X"08",
		X"A6",X"00",X"08",X"DF",X"08",X"97",X"35",X"CE",X"FD",X"BE",X"DF",X"2D",X"08",X"39",X"DE",X"31",
		X"5F",X"96",X"39",X"8B",X"F8",X"C2",X"00",X"E4",X"09",X"50",X"DB",X"35",X"D7",X"35",X"CE",X"FD",
		X"2F",X"DF",X"2D",X"08",X"08",X"01",X"39",X"D6",X"39",X"54",X"C4",X"07",X"CA",X"60",X"D7",X"32",
		X"C6",X"FF",X"C9",X"00",X"C9",X"00",X"20",X"E4",X"96",X"39",X"47",X"25",X"13",X"CE",X"00",X"00",
		X"DF",X"60",X"DF",X"62",X"DF",X"64",X"DF",X"66",X"08",X"CE",X"FC",X"A9",X"FF",X"00",X"2D",X"39",
		X"85",X"02",X"26",X"0C",X"C6",X"5F",X"D7",X"32",X"CE",X"FE",X"15",X"DF",X"2D",X"7E",X"FC",X"80",
		X"FE",X"00",X"08",X"20",X"F6",X"5F",X"96",X"39",X"8B",X"AE",X"C2",X"00",X"D4",X"68",X"DE",X"08",
		X"A6",X"00",X"08",X"DF",X"08",X"10",X"97",X"35",X"CE",X"FD",X"2F",X"FF",X"00",X"2D",X"39",X"C6",
		X"60",X"D7",X"32",X"DE",X"08",X"E6",X"00",X"D7",X"37",X"08",X"DF",X"08",X"D6",X"39",X"54",X"24",
		X"18",X"CE",X"FE",X"73",X"DF",X"2D",X"39",X"5F",X"96",X"38",X"47",X"C2",X"00",X"DE",X"31",X"E4",
		X"00",X"1B",X"A7",X"00",X"7C",X"00",X"32",X"A6",X"00",X"CE",X"FE",X"5F",X"DF",X"2D",X"39",X"78",
		X"00",X"37",X"25",X"13",X"27",X"06",X"7C",X"00",X"32",X"7E",X"FC",X"7E",X"BD",X"FD",X"15",X"6D",
		X"00",X"01",X"39",X"7A",X"00",X"32",X"08",X"A6",X"00",X"DE",X"08",X"A6",X"00",X"08",X"DF",X"08",
		X"97",X"38",X"CE",X"FE",X"47",X"DF",X"2D",X"39",X"00",X"00",X"55",X"55",X"AA",X"55",X"5A",X"5A",
		X"96",X"69",X"66",X"66",X"CC",X"33",X"3C",X"3C",X"0F",X"F0",X"10",X"FF",X"02",X"02",X"02",X"02",
		X"02",X"02",X"02",X"02",X"2F",X"2F",X"50",X"10",X"80",X"FE",X"2F",X"10",X"40",X"FE",X"2F",X"10",
		X"A0",X"00",X"FE",X"2F",X"10",X"50",X"00",X"FE",X"2F",X"10",X"28",X"00",X"FE",X"2F",X"10",X"14",
		X"00",X"FE",X"2F",X"10",X"0A",X"00",X"FE",X"2F",X"10",X"05",X"00",X"FE",X"2F",X"10",X"02",X"00",
		X"2F",X"10",X"01",X"00",X"2F",X"70",X"C3",X"00",X"01",X"00",X"FF",X"00",X"FF",X"00",X"01",X"80",
		X"3C",X"2E",X"00",X"F0",X"20",X"00",X"9C",X"20",X"50",X"6C",X"EC",X"20",X"40",X"63",X"E8",X"80",
		X"1C",X"70",X"F4",X"0D",X"20",X"0C",X"30",X"40",X"00",X"02",X"FF",X"00",X"FE",X"FE",X"80",X"30",
		X"63",X"05",X"2F",X"E0",X"67",X"F2",X"80",X"30",X"02",X"FE",X"00",X"FE",X"FE",X"00",X"02",X"FE",
		X"00",X"FE",X"FE",X"00",X"02",X"FE",X"00",X"FE",X"FE",X"00",X"06",X"FD",X"3F",X"00",X"FB",X"31",
		X"00",X"00",X"02",X"80",X"31",X"20",X"06",X"60",X"DE",X"70",X"D7",X"0D",X"40",X"F0",X"FF",X"12",
		X"08",X"A8",X"18",X"01",X"08",X"04",X"A8",X"18",X"01",X"10",X"04",X"20",X"F8",X"FF",X"20",X"10",
		X"F0",X"10",X"01",X"01",X"86",X"03",X"8D",X"02",X"86",X"04",X"CE",X"D9",X"39",X"DF",X"00",X"16",
		X"48",X"48",X"1B",X"CE",X"FF",X"2B",X"BD",X"F7",X"FA",X"7E",X"F4",X"CA",X"FE",X"9A",X"FE",X"E0",
		X"FE",X"9A",X"FE",X"F0",X"FE",X"F3",X"FE",X"FF",X"FE",X"F3",X"FF",X"24",X"5F",X"D7",X"0D",X"48",
		X"48",X"8B",X"5C",X"C9",X"FF",X"D7",X"0A",X"97",X"0B",X"DE",X"0A",X"EE",X"00",X"DF",X"08",X"DE",
		X"0A",X"EE",X"02",X"E6",X"00",X"D7",X"0C",X"08",X"DF",X"0A",X"CE",X"FE",X"88",X"DF",X"0E",X"7E",
		X"FA",X"BE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F7",X"A9",X"F0",X"01",X"F8",X"08",X"F0",X"01");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
