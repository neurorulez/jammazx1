-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0A4193FDDB0DF08ACAECA7F645CD6330CA553D9FD30F18B3F7E4CC134F6C5DFD";
    attribute INIT_01 of inst : label is "148F6F1DF28145E5D5F3CB20FFFF3CD78FC6ACFFFC95E4DCF2DACEFCA79FCFCC";
    attribute INIT_02 of inst : label is "F480BA3BC3E2F41EACA174D5AF2B4D7B0BCA514BF8BF428D4FCFDCAEECA2C1B9";
    attribute INIT_03 of inst : label is "CA539E39095AA5612FEE05BFFFF7CF70CF2CF2EDE28AF240B9FC07BDCB1FE2E9";
    attribute INIT_04 of inst : label is "BDFABD7E2F5CF38E0E30C0E2F465589787B5E3F4255BB0ACA53B8E14B7CFB3CA";
    attribute INIT_05 of inst : label is "B9947E2CFC71FCA478CB977CA1FED2C7973DFD7E5EAF7F8BDFABD7E2F5EAF7F8";
    attribute INIT_06 of inst : label is "4F352F507C5EC300E06E3CD062431E17E3CD17CA5C7F8BE457CE5C7F8F144D73";
    attribute INIT_07 of inst : label is "F830FFBE0D1461F83CE53AFD5743C6FECAD3847C3C3447C8FFF2FC8FE4F1DBB7";
    attribute INIT_08 of inst : label is "47B28C354EBF57811D11E4F4D077BF439710E7EE0F565A19E788FCDF8005C3FE";
    attribute INIT_09 of inst : label is "C6CA3F3CEC1BFDD7130BD750E60F666365EFAFD5ECE3387A38FA3F3AC05F01C4";
    attribute INIT_0A of inst : label is "FE8EF38C282855707EAFABF852CFEC38F2F4C39543FB83F3D7E2D3BC3A854587";
    attribute INIT_0B of inst : label is "ED69453C9C374B7D7A3DF7EF0E1795876BF5ABF7DAE8EEFCA7C72DA6C33DBC38";
    attribute INIT_0C of inst : label is "EDFD7EFD5BDF16D7FCFCB3FFFFCF30B2E9F11DD5169555692D55669555485C17";
    attribute INIT_0D of inst : label is "05FB0BB429EAB44D411152347F73CF1D3DC0F0CB3C71C70C33FF14552CBCD7C6";
    attribute INIT_0E of inst : label is "73826134D07CA29C9E171D3FBFC1F0F739CA0C270E99555695556955548E171F";
    attribute INIT_0F of inst : label is "3DECF4D7E4FB3F5C3CFD70CF7221FD8A17C55BB87D735144175EB64FF33F2BF8";
    attribute INIT_10 of inst : label is "FE475B1E6C4569861B65B69848FF23FD4C101CCFD6AC503ADC2C3FF471055F9F";
    attribute INIT_11 of inst : label is "B1E8833F75B1E6C6D645D464C60CFD75B32C79B1B5761CFDD6CCB1E6C6D7F60C";
    attribute INIT_12 of inst : label is "CF8EFF69079833DC3E4D9833DD5C873FFD4B57EB833F5D2CDB1E6C6DF65756CC";
    attribute INIT_13 of inst : label is "57DB77ADD1CB6703EB556034FCD3F97E3CF5DBCD0E4F7D938FC363CFF396D594";
    attribute INIT_14 of inst : label is "D7EEE8EFA23CFF537DAB3FC3D67B0EBC39556626EE6AA22AA15774057DDDDDE4";
    attribute INIT_15 of inst : label is "F7F7FBF7FFFFFFE7EFE3E7E3EBE7E3EFEFEBE3E7E3E875DD8F3FD155FEB0F729";
    attribute INIT_16 of inst : label is "FDFFCF3690DD5503D03527544D55555445544DE53355515455113007E3F7E3FB";
    attribute INIT_17 of inst : label is "BFFAFFBFFBC1E50775144B1FBFFBFEBFEBFCBFDFFCFEFBFFBFFFFEFFEFFDFFCB";
    attribute INIT_18 of inst : label is "FF7CFBFFFCF7DF17945D545513C76FF6FF2FF6FFAFFBFFBFB6FF6FF7FF7FF3FF";
    attribute INIT_19 of inst : label is "7EF3EFFEF3CFFEF3EF7CF7FF7FF3EFFDFBFF7DFBFFFDFBEFFDF3EFFDFBFF7EFF";
    attribute INIT_1A of inst : label is "FFFDFFCFFFFFDFFCFFFF07941D5590D146F9EFBEF9EFBFFFFBCFFEF3EF7CF3EF";
    attribute INIT_1B of inst : label is "7FFBFFBFF7FFBFFFFF3FF3FFFFF3FF3CFFFFFCFFCFFFFFCFFDFFCFFFFFDFFCFF";
    attribute INIT_1C of inst : label is "1D149C51555517945E5965955357575111540471796507555957755551047BFF";
    attribute INIT_1D of inst : label is "D552594DE595516511051555145574507955925940D555557765D51440451455";
    attribute INIT_1E of inst : label is "55DCDE5545555C5D551FD5155474537955555379659651D44D04591455D1D14E";
    attribute INIT_1F of inst : label is "C1E52756554DE55555541C9E517975957555507079941E5975445D5517955114";
    attribute INIT_20 of inst : label is "59D45759455517FDBFFFFDFFFFFEFFCF7795DDD515D074251055474F9554155D";
    attribute INIT_21 of inst : label is "455136F925551D4565D4540D4E595547795556554555D5D457595554D4575575";
    attribute INIT_22 of inst : label is "06EF83B7CF3405867A79A3154FEBDDD7735645541DE5555111767D6557964940";
    attribute INIT_23 of inst : label is "4D443EEA1504C501FB9AB04D051D2B04D445A141555B11BE1CEF5EF05F3C13EF";
    attribute INIT_24 of inst : label is "F5FFE0FF0644797A5EFF2E847EEA1407EEA144FBA8517EEA554457EEA141FBA9";
    attribute INIT_25 of inst : label is "FFC3CAC3694D815D8744615D175B47F75D7828B33CCE33CCE338CC307459C1DF";
    attribute INIT_26 of inst : label is "7D9FD2A247F7343DC1FFFBBD725E5F0EFBB4F56C1FCF07F7C17DF47FFD1FDF07";
    attribute INIT_27 of inst : label is "501A45FFFFF05A51704555A151C4C456AAAA6A5441555B57D163F09EEBC21DF3";
    attribute INIT_28 of inst : label is "7061F0DFA6DDC17F5F8FC33F0DFC0F7E0FDA5571501AB5575536A56B5A51355C";
    attribute INIT_29 of inst : label is "D472457FE9B5C56A6FFD5AB2ADAB2ADAB6ADA994D441B578D1FDCEDF5C37E5B7";
    attribute INIT_2A of inst : label is "B76C10E3FEB86AE29955D416D5E347F7D17F78F47F78F0FFF702FF8374709397";
    attribute INIT_2B of inst : label is "4597C1DF1F65D1FCF05F7C13FF06EF83F578B2CFDD5E38BE2BCAC1304FEC137E";
    attribute INIT_2C of inst : label is "7D1FDF0E14B1CF8F2CFCBAEC3F8AA25E6ACF33C3EAE9EF8F6CB7FCF6CB8391EA";
    attribute INIT_2D of inst : label is "6A51D9405761C51AA5D456AD45C04D2B151D45A557515B579580A67A9165F47F";
    attribute INIT_2E of inst : label is "F6CB8391EA4597C1DF1F65D1FCF05F3C13EF06EF83B578FCB2FC6840D45EC744";
    attribute INIT_2F of inst : label is "507117B1D11AA5D446AD44D051D2B151D44A557511B57CEA2ECAF9EF8F6CB7FC";
    attribute INIT_30 of inst : label is "1D1691F245C5D3FEB13C13C199789858FD97BFD3F47F7C1FAF05E7C13AE0ADA4";
    attribute INIT_31 of inst : label is "5AA152A856A81AAC453FFFEC451AAB51555747FA140750417F6A5575016FFD5F";
    attribute INIT_32 of inst : label is "54CC6468C1F70C0F7175B7F3C7AFA5BDA543AA45FAA153AA15FAA0FF6A555AA4";
    attribute INIT_33 of inst : label is "E3BB197E3FEC38F3FCFFBC62CF8F4B3C72A4ACF18B3B0B2B577A6D7DDD39DE49";
    attribute INIT_34 of inst : label is "B179D0BC1B9F8D3D0F3E3FB32ACC2F0A83BE6A8979F4F0F2FF0B2CED3AC387E0";
    attribute INIT_35 of inst : label is "E8453B1EA114EA042A8106ED0FEEC8E5E51FA8EA3BC3CB1F2F4EC2B8159C1F9F";
    attribute INIT_36 of inst : label is "B0B8AE28A7E87AE704EF4E1E3DFBBB0704EBD12F68ED1C02FEC29B8BE3E8F3F4";
    attribute INIT_37 of inst : label is "63FD2CE7F3F2B43FAEC6CFEE306E7BCAD0FB4EBC452854C56AF114A11D5582FB";
    attribute INIT_38 of inst : label is "57E930C754FA455D5704566E28AF07D8FF6B39FCE4E07B43FAEC6CFEC13AF8D3";
    attribute INIT_39 of inst : label is "1FF654BED3DBA55C15BBF9BED45A45156FBF9B1C106AA154D35405D0DAB55D14";
    attribute INIT_3A of inst : label is "E2F93E40BCEF9EFAE7BFB0ABE4E7F719D3E9B70A86C9503141F107FFC68DA45B";
    attribute INIT_3B of inst : label is "66913EAB420080226FFE6F95FFF3BB3BA5CC792FD04ABE2CEBEFBEFA6AFEA0F8";
    attribute INIT_3C of inst : label is "C837912B660B20AE1F2883A8ACE2C56EBCBBDBE8D1777F3BDEFDF0E8DA7B9DBA";
    attribute INIT_3D of inst : label is "8F7BC2978288FEEC2BD3FBC3FFF83D2E0F0B720F4CA5EE4E40EA4ED52A683CEE";
    attribute INIT_3E of inst : label is "C21C178C2B05B7835647668A2BA87F06E3FFAB8F9EF3A2F8FC3A8EB83E3BF0AB";
    attribute INIT_3F of inst : label is "D54E8BFDE8FE3FB12C8F5E661D39194CF6CCFF166E328F13F060D5E9F0CFC3F8";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "CDF442AA237EBA47BCBB86902851863AB0DDB258388753415D4EC9E3A53C71C0";
    attribute INIT_01 of inst : label is "2F56388DEE31C7170DF33DC3B6C9ED7F3EE5ACCAA85FA888AAEBAC7B8B5A8A8D";
    attribute INIT_02 of inst : label is "BB4339F23D1E0E9CFB8DD2673EE1267337B8DDFCE72B2F0B78083D6BE8F68F07";
    attribute INIT_03 of inst : label is "B8BF1DD1EA6AA64AE0FC2732CB2CB20EF0E2CD0A9E7C8FBF8583A7337FD8CF20";
    attribute INIT_04 of inst : label is "7FB17EB9DFAF8E7AFBE3BFBCA75E72A73DB9C999AA70F13B8BF274DFC61FF39B";
    attribute INIT_05 of inst : label is "FB1871C3425DBB07BF7C5C7BC1CCBDB3DC58FFF9FE5FEE77FB57EB9DFAF5FEE7";
    attribute INIT_06 of inst : label is "BAAB92BDEBDFBEFADABCBBF45603FBEBCBBFD7BC70733CC777B870733877D5C7";
    attribute INIT_07 of inst : label is "486B82521EDF536C1ACCF1F7158E04BC8F8E07E7677BF6B380AC2B38C7BE779E";
    attribute INIT_08 of inst : label is "F181FACF3CFFF1C31FBC2FE7ACFF7FF5539D5323D5F4D353C9051B91887DAE09";
    attribute INIT_09 of inst : label is "BCF0E0F3CFE3E7D191FFFD3DFF8BCFBDECF83FFCFC0AADA747C1FAFBC3DB01CE";
    attribute INIT_0A of inst : label is "CA74FDB852D35D7FCB02C0B2DFF9BCF3BC7ECD1D7B32FB0F6B9D67FCF29D41BE";
    attribute INIT_0B of inst : label is "B76B47EBBFF57BE7FDEE9BEF3CFD5C4D17DCC7D72C9CBABB8ECDFF9DC1EFFCF3";
    attribute INIT_0C of inst : label is "DD61E1F742B8FEBB9463ECB28A2B038C1586ACDE06AFFFEAA6952285556B7FEB";
    attribute INIT_0D of inst : label is "FAE9FC68E95F55848617A2FBFE5EFBCE28E2B4DF79E3CF2CB3FF0377E3017E3F";
    attribute INIT_0E of inst : label is "9FB2AAEBAEF39E38BBEBB7B33C8BE3EED3B8820D8EBAFFFEA555285556BBEBB7";
    attribute INIT_0F of inst : label is "583B361CC631F777B7DD5ED600884049B903DE255DCC57041C71A270060B0092";
    attribute INIT_10 of inst : label is "CB7E69D8A7FDFEFBECBEDBEEB4CA3BAB8C1208A430F57357F8CC5A18C9B7DC5C";
    attribute INIT_11 of inst : label is "9F747B32E69D8A7F27759FFA8DECC9E69EA7629FC965ECCB9A7A9D8A7F2725EC";
    attribute INIT_12 of inst : label is "FC7CB27DD817B319F09017B31B487B32AB9C95B07B3279A7A9D8A7F207A23278";
    attribute INIT_13 of inst : label is "66E7BA5CCD208382A17D73D3E70FDEB1CCA48709EF7E7A5E0C9A9CCCAE3F248E";
    attribute INIT_14 of inst : label is "BCDCF4BE51CCCAF2AB6F32AE196F34BCD1DD37B7EA3EA73EADF67B666AEAAA16";
    attribute INIT_15 of inst : label is "9293DF9F9BD79FA3A3E3ABABAFABA3A3ABB7BFA2A3E3219973329DDDCC8CA22F";
    attribute INIT_16 of inst : label is "FFBFFBAD36B69D19BEFE9DF6CEFFEFFFEEEEAF4DA3BFFBDEEBAD3087E3DFAAD2";
    attribute INIT_17 of inst : label is "EFB7FFEFF6E70C9DE7B42FACFEDBEDBEDBFF7FFBFFBDC7ED7FCBFDBFDBFFBEFF";
    attribute INIT_18 of inst : label is "BBEFBACBEEB2EBCC33338EECCFEBFFBEFB6FB2FF5FFEFF6F7DFBDFFEFF2FF6FF";
    attribute INIT_19 of inst : label is "EFB6FAEFB69AEFB6FBEDBEFAE9A6BAE9AEBAE9AEBAE9AEBAE9A6BAE9AEBAE9AE";
    attribute INIT_1A of inst : label is "CFFBFFBFF8FFBFFBFF8FEC33B38C0DFBABE9A69BEDBEFAEBA69AEFB6FBEDB6FB";
    attribute INIT_1B of inst : label is "7FF7FF3FF7FF7FB3FB7FB3FB3FB7FB3EFEFFEDFEEFEFFEDFFFFFFFFCFFFFFFFF";
    attribute INIT_1C of inst : label is "EFFAF6EBFDBFAC3274E3CF357CBDFDFEABA2EAB9E38E8DBFF355DFFBFBBBB3FF";
    attribute INIT_1D of inst : label is "7DFDF7EB4D7BFFC7EFEBABFFBBFEBFE9C33D3CE3A07DBAFBEBFDFC1FFFEFEAEF";
    attribute INIT_1E of inst : label is "EFFE34DDEEBBEE6EFF977FBBFEBFEBC31E7DFAD79F7CD98FF6BEFBAEEFFAFFA0";
    attribute INIT_1F of inst : label is "E70CA9BCEF6F4DEFF98EAE70CBD39F357FFA3AB8F13E34D7FFD6AE7FAD35FDAE";
    attribute INIT_20 of inst : label is "9B7EF8F367FBBFCFBECFEFBFDBFDBFDB4C31379DC7FAB4AFBABBCF673BFAAEFF";
    attribute INIT_21 of inst : label is "4B3FF703CEF1737F8C0FEBFDF6F3BDE4D3FFF8D9EFBED37EF8F37F9A7EF8FF7F";
    attribute INIT_22 of inst : label is "FACD4DDF88F36D14E3E38118C0F94FFB44F0FBBBDF0CFB3FFFB4CF8C6D34F3AE";
    attribute INIT_23 of inst : label is "44D5146A0B545904558AA45551D66A4554C5A0D287682571786C8FBF9D5FEB57";
    attribute INIT_24 of inst : label is "09FBF1B32BA571C58FAE6E9F576A295146A19851A8D1D56A4904A156A38551AB";
    attribute INIT_25 of inst : label is "CDCE3CBCEBD79635997DEDCC9C73BEC1D5833C7A0286B16C7A1282B132739DBC";
    attribute INIT_26 of inst : label is "8FF06A99990AA99BFF4659AA789C73F76D5BF9CFE707F8C5FE737B9C1EFB07FA";
    attribute INIT_27 of inst : label is "115A4755555C5AD1DDD30DA7504544FEA1412AAD44CA296DC9C0DD2B73743630";
    attribute INIT_28 of inst : label is "7F537F66EA55FF519E376CFDB3F6F5FD367AD6D7315A9D6D7156A0A9AA6615B5";
    attribute INIT_29 of inst : label is "960A27FF2B9A5A2AE5569A91A7695A7699A66BB44D5296C3EFB07D9ADFD9B695";
    attribute INIT_2A of inst : label is "55EFDDF5A291EA46BA1C785A5B0FBEC14D8D90D39DD0DFFFF5F0FF4D5FF07BF1";
    attribute INIT_2B of inst : label is "271C9DBAF7C7EFF07F9C5FEB17FACD4CDD07FE7835B0EF2BC23CCFEF7CCFD59F";
    attribute INIT_2C of inst : label is "DEFB073DF70F3C74D2C3C8945F26999C97C3AE0E05100F4B0740BCB875CAE9CF";
    attribute INIT_2D of inst : label is "AAE17AB1C9665DFAAA7472AB4755466A136747A871D1E96D678EEA72C9C73BFC";
    attribute INIT_2E of inst : label is "B875CAE9CF271C9DBAF7C7EFB37F9C5FEB07FACD4C9D0783FE63E8557475597D";
    attribute INIT_2F of inst : label is "455265565F6AAA5982A998551D66A136598A87166296E319DB85200F4B0740BC";
    attribute INIT_30 of inst : label is "EC9C7F75F9D7103E17ACBAEAA872A870601367903BEC1FF767F9DDFEB45367A7";
    attribute INIT_31 of inst : label is "9AA732A91EA96A8477555554774AAA573F3D455A2951504555EA871A54AFE5B8";
    attribute INIT_32 of inst : label is "2BB16F2BFEB73BF44F9779DE8DC98DBBAC95AA895AA731AA475AA555AABB8AA8";
    attribute INIT_33 of inst : label is "9F3EF1CDDABCF3B1B3BABB8F3856370E112CBCAE3C3F34C1E7C0F5F02059D8F0";
    attribute INIT_34 of inst : label is "F272733FEB16F9CCFCD1D02AC073CF300C6A1A6670B893BFEF3FEFC9CBCB3C23";
    attribute INIT_35 of inst : label is "28775125A1DD5A452A811EDFFCC947C716F32789F23C30493F6D82FBA73FE716";
    attribute INIT_36 of inst : label is "F34749E7CD1280CFFAC9F9DBDB47C20FFAC19FC0678CCA3C0F8D3E3DBE47FB27";
    attribute INIT_37 of inst : label is "1D2CBB45BCEC3FF21939F4CBFFAD53B0CFC67294776B54546A51DDA125D0BC32";
    attribute INIT_38 of inst : label is "A16A554D7D5A4846E144BE5CE788F8074B3ED16FF23A73FF21939F44FEB76F9C";
    attribute INIT_39 of inst : label is "FCADAE7FEBB0A7451D995F95747A5B686595F955146AA474658D3A514AA7456D";
    attribute INIT_3A of inst : label is "8189AB23FB4EB28B24A3E24B22CDAEB3AF2B12244A88C8FDDE191F002BBE8738";
    attribute INIT_3B of inst : label is "2C38A8F0D1E058023EF26886ABAB262718CD2C9FA3ACBACB48248283AACB6286";
    attribute INIT_3C of inst : label is "4458C995067C0BCCEE926C07FB480D5C9849872BAF22E8A228A0F2BC9A20890A";
    attribute INIT_3D of inst : label is "B37BC933CA16CCBC3EEF9EFFAAA3AEF8EBFE2107EA4FE9EBEE9B2BA99E95BD9F";
    attribute INIT_3E of inst : label is "44243FEC937F28C3FE31EE79D2F2CBACECBC73B3A4FE6FEFBCF27438A1A1E263";
    attribute INIT_3F of inst : label is "7FC2B6ABB0BC28E3DE5DDF953558F3E9C9ECCA3DE503FE3EA0117E92C3AA8FBE";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "67CBF87BEB1FED2E3AA321421A7D37733214D1B65569FAC3DF1DDE768D85FBE4";
    attribute INIT_01 of inst : label is "97EC3D638E90DFEFC5559F4160E0D1D3574531F555111A3307123223A601E1EC";
    attribute INIT_02 of inst : label is "1F6B8E799DAD9C7EA36417EFB8C97EF9D6320476B53E1D8D11E1D6BEFEEB669B";
    attribute INIT_03 of inst : label is "32578FF856155A09C9661FB8638E186F3EDB2D8D679E65D76B671F9B3C766F98";
    attribute INIT_04 of inst : label is "D7CBD58E7571E7DD5C79C557F5BAF96F947BE47A59FB9A632579FE47ADAD9BE6";
    attribute INIT_05 of inst : label is "7DF4FACBE584E3A126FEBE23E3E6C6DA7EB0F7C7F1F5E39D7CFD58E7570F5E39";
    attribute INIT_06 of inst : label is "D0CC4BF25D29451F073E170CEE814573E170423EF8F9BE611236F8F9B6916FE2";
    attribute INIT_07 of inst : label is "BE1DCFAFA45552581320F9F416CFAF6E061F95511191551FE54751FE6546D752";
    attribute INIT_08 of inst : label is "C3D77D143E7D118930F0B7E3D097F55B41C6D10A5727BEFEFBC355389015773E";
    attribute INIT_09 of inst : label is "163AF9FB6D7C541665876105954FA77B4061DF446A70CEDFAFE3F8F9A946231B";
    attribute INIT_0A of inst : label is "E39E5632CDF9101131DCF71C0C39E67B0D5B6F811C995C9E50FD50E678263411";
    attribute INIT_0B of inst : label is "D4422251CD595DF74755D4199E43504927D067959EE6A3A32F01E4FD05E4E679";
    attribute INIT_0C of inst : label is "D6C519F44DCE45DCD4F97A2863BC36F8EB4EA400400000A245404A0000914D78";
    attribute INIT_0D of inst : label is "5E15769903D7B31D3CD92075E3D5144F80EBC8CBA849A69A68AA0914EB27D391";
    attribute INIT_0E of inst : label is "D518CC000145E5B2057454E99A25197CFB32CBACC010000A2FFFA00009157457";
    attribute INIT_0F of inst : label is "B07F0DB66FBA3DF748F7DD2C1155D52B61D044297FF2D781FFDE011DDDB3F73D";
    attribute INIT_10 of inst : label is "F5501541951515C79571E75C45F57456890C73514F3025B732C09734045136B6";
    attribute INIT_11 of inst : label is "546A747D01541953155021D221D1F40154550654C581D1F405515419531789D1";
    attribute INIT_12 of inst : label is "961638B545D747D459A4D747D433747D56AC50E9747D00551541953157180551";
    attribute INIT_13 of inst : label is "FEF9DDC7714D37E57D44D9C45713DC79C15227D4D15F35879F4CDC1F57831422";
    attribute INIT_14 of inst : label is "1176E219A9C1F518C0707D558719B6E6F8149991FF1FF19FF448118FEFFF7FF8";
    attribute INIT_15 of inst : label is "F3FD79F17377FF5F53DBDBD7DFF7FBF3F7D3F5DFD75D8102707D545366F60CF8";
    attribute INIT_16 of inst : label is "DF7DF76F3DB0CC34F87E4B7D7FC3BD3EBF379BCF6F74FFB3FDD52617DB575757";
    attribute INIT_17 of inst : label is "DFFEF7DF7DD30C4EBB78192EBFEFFEFFCFFF7DF7DF7DE7FE7DE7DC7DE7DF7FFB";
    attribute INIT_18 of inst : label is "F5975975D65D77AE3AB7DFFDE8E72FFBFFBFFBFFDF7DF7DF71FF9F71F79F79F7";
    attribute INIT_19 of inst : label is "D65D77D65DF7D65D77DE7DF5D75D65DF79F79F79F5DF7965DF5D65DF79F79E79";
    attribute INIT_1A of inst : label is "77FE7FF7FF7F67F77F773E38F7DDE1CFC7D779F5DE7DF5D679F7D65D77DE5D77";
    attribute INIT_1B of inst : label is "DF79F5DF5DF59FF9FF9FFDFD9FD9FDDD7DE7DE7D57D67D67FE7FF7FF7F67F77F";
    attribute INIT_1C of inst : label is "9F7A8FCF9F5F9D367CC38F3DFF31B7C84FD44878E38D9F7AF3DFBF3F64EA7DF7";
    attribute INIT_1D of inst : label is "DFBFCB67CF32EFCC87C04B28FF7C7DEBD34FB6EB62DFB2EBF1AFF1BA7914ABF5";
    attribute INIT_1E of inst : label is "75FCFCF3F7131C05DF0FFFFD7E7DE2D36CBAF2F30E3CFF52F8D1CEE3FDFDF7A4";
    attribute INIT_1F of inst : label is "CB4D1BBCD7CBCFF5FBD31C34D1F37F3ECD7F6E70D3343CFFFD6C95DD2F3FF3D3";
    attribute INIT_20 of inst : label is "B35DF8E3779B53F6FF7FF6FDCFDFFDEFFC33FAEE8D77BC37FC7F4FFF36FF5F9F";
    attribute INIT_21 of inst : label is "20CBFDF3CC7FBFFB0FFFCE9FB7E39D9FD32EF8D11062F35DF8E379B75DF8E779";
    attribute INIT_22 of inst : label is "57217515C65912FF8EBE3365975550F75F7CFF33D3CFF0F85F3CFF0F5C30DF07";
    attribute INIT_23 of inst : label is "7D667FE849A1E8F1F790292C84CCA292E352056485B3977DD0CEC3F5E15D7467";
    attribute INIT_24 of inst : label is "DE1D9A36525DFBEFC3C884273FE8628FCE8681FBA188BCE8183287EE843CF7A0";
    attribute INIT_25 of inst : label is "114796F5436D327D233644687EFB5D3D4479AEFD97E6D9FE5DBBECDAE1F9E6DE";
    attribute INIT_26 of inst : label is "C1FE357B8E8D9830D4D5BD7DC4BEFB5C5BDF3BED70675E1DD78775719D74F75E";
    attribute INIT_27 of inst : label is "5E90B7FFFFF54888B685A6098DF3D264089D80867068711587EEC79E7B162746";
    attribute INIT_28 of inst : label is "755375E59BD5D43161B9C5F317CC79F1DC50883B1F2038832DB80A0380A0720E";
    attribute INIT_29 of inst : label is "0022313D4134E2C04FFD203E0C83E0E83A0D8107D6671179D74F78401D796AF5";
    attribute INIT_2A of inst : label is "B57D449B343440F0114DC3CC45E75D3D64D19059F11251E7C1196C75D5AA0A53";
    attribute INIT_2B of inst : label is "1FBEE6C45434D74E75D3DD74E7572177113B0E7E545E55FC5B9645513E6D4B9E";
    attribute INIT_2C of inst : label is "1D74F519472F9EBEFBA5E6EE35997BBE4E6CC7A5BBD86661F1F1EA1F8F9797EA";
    attribute INIT_2D of inst : label is "4008D3165788F95032E2240A22F21CA2CC2E22053788B115940698F987EFB5C3";
    attribute INIT_2E of inst : label is "1F8F9797EA1FBEE6C45434D74475D1DD7467572175113BE70E594123E22FE336";
    attribute INIT_2F of inst : label is "12342BF8CD9032E8140A81C84CCA2CC2E810537A071159BE4E2BC86661F1F1EA";
    attribute INIT_30 of inst : label is "787E75C1D72FBE5B887A67A561F961FAC4FCF7FE75D3DD5C775731D5CF5DF503";
    attribute INIT_31 of inst : label is "288B1E228A23203F16FFFFDF16F2228B1B1F37F8628F853CBF405378A3CF7456";
    attribute INIT_32 of inst : label is "82ABFC3DD7C51F7E55317DC7C9EEE45D0D8F8882F88B1F88A2F88CFF80991888";
    attribute INIT_33 of inst : label is "6598FBE940E67B8319CFE36CB2AC3C1538B9E67DBAB9B2C9DCACA73766FB3FBF";
    attribute INIT_34 of inst : label is "9B8E4B8D70F71D565EDAF93CE91959BAC6FF65EEF81E29C7799455ED526EBE41";
    attribute INIT_35 of inst : label is "4316FFCD0C5BD0B66214F43E766EEB6F91F9B9EE599FB201B292EB9E5F8D78E7";
    attribute INIT_36 of inst : label is "9B232679E784EA635C1516456DE1ABA35C1DD4E93966469E96ECB8F96E69CEB5";
    attribute INIT_37 of inst : label is "7D876363458EB9D9AC9F36AC7573DA3A65EB543F16E193E080FC5B8C8C131E9A";
    attribute INIT_38 of inst : label is "87E0BCD706F8323E47B190B679E6767F61F8DAD1A565FB9D9AC9F366D58D71D5";
    attribute INIT_39 of inst : label is "4E019046E38D004E593BFB3DE22809A14FBFB39ED9488921CB5653C4F0204C26";
    attribute INIT_3A of inst : label is "AFE2BE54E3EB28638E08B9A383EC0C78B780CD9A5C2BE4C7D613B15556B03C2D";
    attribute INIT_3B of inst : label is "03FE416D0BBACCBCDD780E0B5555BBBD966EB966647AA7A3E18E082C40E19BAB";
    attribute INIT_3C of inst : label is "64978440A03627655869DC8D63E6A1FA01D22F81B480017C5F04212AC03D0CD0";
    attribute INIT_3D of inst : label is "1716668AEC8FA66EB837F837C006C35DB0D7CD26F1A0FF5ED5FE5EE5599D7A1F";
    attribute INIT_3E of inst : label is "E13E807668D0D54156D0F29E5BB9619645F7D917DE57BE5B967B96EECACABBF9";
    attribute INIT_3F of inst : label is "41080C006A188388706D095525B06833FD81F545D5382E7156504306E9A065C7";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "7AD19EAD5E5DACFE76A727F6634127207E55E0EA58B123044436C972E3888AA4";
    attribute INIT_01 of inst : label is "749AFDC99C80CBFBD022DB79AEBBF8835E82ABBF3FD5B7BBAEBA72A726CABAB9";
    attribute INIT_02 of inst : label is "E41FAA6F5EBF932AE7E0289AA9CA89AA9A76503E297ACF9D4ABA82FAB9AB9CAB";
    attribute INIT_03 of inst : label is "72DF9EC93D3FF170C9ABCAAEBAEFAEBFBAFB6CA8A69BD653EEE4CAACFE2EBFBF";
    attribute INIT_04 of inst : label is "EAAEEA287A8886584969A4A7ED29ABDA80C6ACE6F7ABA6A72DFAB2036AAEA6EE";
    attribute INIT_05 of inst : label is "EDB0ABFBA720A7A42CBAE227A2AB87C6E26B3BAAAABAEA1EBAEEB287ACBBAAA1";
    attribute INIT_06 of inst : label is "9AEDFB766C1BB6DCA3DBDA95F1960A7DBDA9027A88AAFAB4027E88AAFE940A26";
    attribute INIT_07 of inst : label is "B9A53EAE685424A96763EAE9D26FA3AB6A7FB425A5A1425BE696A5BEB4A58AA2";
    attribute INIT_08 of inst : label is "93E2BA60FABA5F940964B7E7A527AA428CD1AE1869410524D3796916038094FA";
    attribute INIT_09 of inst : label is "58BAF9EBAE62E958999BB210B2DC36E223A6AE97A9A2EAFA9BA2FAFA940A5095";
    attribute INIT_0A of inst : label is "BA9FC7870BC800792DAB2ACB4CB2E9FB6DBC9E954DAE5D9CA6EDA6A9FA800182";
    attribute INIT_0B of inst : label is "E96800258E767A8A2AFA28AA7E068392FBA7BAA6FBA9A6E76A92C9AB96D9E9F8";
    attribute INIT_0C of inst : label is "B8A83EE97ACD56EAD8B5F3BEFBF6327BF3EF9D01069555696400669555580E6A";
    attribute INIT_0D of inst : label is "9ABA3AE76855500400000639BB629A7DEBDF649E38E3CF2CB2FF5400CBE58356";
    attribute INIT_0E of inst : label is "A3DEEF6DB7A4A6C7896AE9CAF9BEBDB1E876FBE3FA9955569555695555896AEB";
    attribute INIT_0F of inst : label is "6B7F6BAEFABC6AAB61AAAD9AD3B99573894152CB0E3CCFE3EFBFA40A926E6ACB";
    attribute INIT_10 of inst : label is "BE563A5B690020A28A20824A0BB3EEFC688E3B29454AB02AD7D96BE009802AEA";
    attribute INIT_11 of inst : label is "A4A3B6EF63A5B692C252A3EFB6DBBD63A6E96DA4B0AACBBD8E9BA5B692C2EADB";
    attribute INIT_12 of inst : label is "BAFAAEB96E8B6EDEEB6B8B6EDD3BB2EFFC6B03E5B6EF58E9BA5B692CA2CA8E9B";
    attribute INIT_13 of inst : label is "9BDF77BDD07AEE6CEE5534D9EB26AB2EDBF2AAFCDA5B4FDEBBEEEDBBFE82C2A0";
    attribute INIT_14 of inst : label is "41ABE3AB8EDBBF5EE9A2EFFE8A2A7AA9E9552266EE6AA22EE00AA1B9B9D999EB";
    attribute INIT_15 of inst : label is "A6A2A2AEAEAEAAB6B2FAFEBABAB6BEBABEBEBAA2AAA8A8AAB6EFD002AB97AEF8";
    attribute INIT_16 of inst : label is "ABAAB8EE3BBB9FFEFFCFFEFBABEFBEFBFFFFFF8EFAFBEFFFFFF0A286FAEABAAA";
    attribute INIT_17 of inst : label is "2AA2AA2AA2338ECEF7FFF3FAAAAAABAAAABBAABAABAAAAAAAAAAAAAABAABAABA";
    attribute INIT_18 of inst : label is "AA28A69A2AAEA8EE3BBBDFFFBEFEEAAAAAAAAAAE2AA2AA2AAEAAAAAEAAAAAAAA";
    attribute INIT_19 of inst : label is "2CBAEBACBAEBACBAEB2EBAEA28AEBAA9A69AA9A69AA9A6BAA9AEBAA9A69AABAA";
    attribute INIT_1A of inst : label is "9ABBAB8AB9ABBAB8AB98EE3BBBDFFEFFFFAAA2AA28A2AB2EB2EBACBAEB2EBAEB";
    attribute INIT_1B of inst : label is "AAAEAAEAAAAAEAAAAAAAAAAAAAAAAAAAAA8AAAAAAAA8AAAABBAB8AB9ABBAB8AB";
    attribute INIT_1C of inst : label is "F3FFBBEFBEF7EE3BB861863BFFFFFFFFFFFFFFCFE38EFEFBE3BFFFFFFFFFEEAA";
    attribute INIT_1D of inst : label is "BEF8E3B38E3BEFAFFFFFFFFFFFFFCFFDE3BE1861B7BEFBEFBFCEFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFF3B8EFFFFFF3BBEFE2FBFFFFCFFFE3BEFBEFE38E38EFFFF7FFF7FFFF7F3FF2";
    attribute INIT_1F of inst : label is "338ECEF8EFB38EFF3FFFF378ECE18E3BFFFFFFCDE33B78E38FFF7BFEDE3BEFFF";
    attribute INIT_20 of inst : label is "FBBED8E3BDFFFEA8AA9EB8EA9AA8AAA8FE3BFBDFFEFFCFEFBFFFECF61BEFFFFB";
    attribute INIT_21 of inst : label is "FFFFCCE382FB3BEF8EFF3FF339E1BEFDE1B6D8EFFFFF37BED8E38FF7BED8EF9F";
    attribute INIT_22 of inst : label is "98AEB626CD65614535345F16CFA2A93CFEF82F9FFF8EEBFFFDCCEB8EFE38E3BF";
    attribute INIT_23 of inst : label is "0400155A00004000555A9004000429004000A000001ACFAF88ABDAF98A2E6A8B";
    attribute INIT_24 of inst : label is "9CAFA6BEC6CFAA2EDAE9AE80155A000155A000556800155A00000155A0005568";
    attribute INIT_25 of inst : label is "A6C61BB5680580058100601B22AB9BA65A2569B37CDD374DF27899262CA896DF";
    attribute INIT_26 of inst : label is "AAE29FF768A66668E5EABEFEAF628B9EABA986AE668B98A6E6A8B98A6E6E9B99";
    attribute INIT_27 of inst : label is "000A005555500A00100000A000404006A5556A0000001A80B2AFF7FE2FDF4AAB";
    attribute INIT_28 of inst : label is "7926B9CAB6D9E576AAF2D6EB5BAD72AADD9A0010001A90010016A0290A001004";
    attribute INIT_29 of inst : label is "88D1F56E6990406A65541A91A4691A4691A469804001A825E6E99B8A0E72A1B6";
    attribute INIT_2A of inst : label is "362E50B696946A5298004006A0979BA6F48BEDBD8BADBDAAA7D7AAB7A465C6C2";
    attribute INIT_2B of inst : label is "CAA296C96660E6EDB99B6E6ADB98AEB765EF6DBE5A0969F97E1BC5213ABE5B2E";
    attribute INIT_2C of inst : label is "2E6E9B1D57AEBEFADB27AFA962FFF762FA9C1FBFA6AFBE1E6DADA9E6CAB3B2AE";
    attribute INIT_2D of inst : label is "6A0058000160401A904006A400400429000400A001001A8340B5B7AAB2A8B9BB";
    attribute INIT_2E of inst : label is "E6CAB3B2AECAA296C96660E6ACB99B6E6ACB98AEB725EFE76DB5680040054100";
    attribute INIT_2F of inst : label is "00100150401A904006A4004000429000400A001001A8352A7E76AFFE1E6DADAD";
    attribute INIT_30 of inst : label is "4B2AA7AA9EA8AA6AC82A02A3DFABDFA8ABAE9BEA79BA6E6ABB9AA6E6A8AD89A0";
    attribute INIT_31 of inst : label is "0AA002A802A81A9400155554001AA9000001015A00010000156A0010006AAA0D";
    attribute INIT_32 of inst : label is "9598D92CE6631B7A5060A2F7D2BAF5FDA001AA005AA001AA005AA0556A000AA0";
    attribute INIT_33 of inst : label is "A6F9FA2D7AA9FB62AFEFA7ACB6DAF616099CA9FEB2FA7EEAC23414D333209935";
    attribute INIT_34 of inst : label is "A6A99FAE6E9BDB597EEBE9A1EA5D4A7E94A2FFDD8BE7BFEEBA7AEBEB5E9CBE6D";
    attribute INIT_35 of inst : label is "68001505A0005A002A80062D7ABA9FA8A8FAE9BA6F5EBABCFA8E9EAE3A8E628B";
    attribute INIT_36 of inst : label is "A7EFEA69B8BA2DB39BA64A4A5E2EAE739BA6B5F969B979CF9E9FA9B2AD9FECAD";
    attribute INIT_37 of inst : label is "6CB9A726A69EB5EBFEDAB2BF79BBEA7A97EED694002800406A5000A004018FAC";
    attribute INIT_38 of inst : label is "01681041005A00040100062B29BD7A4B2E69C8A9ACECAB5EBFEDAB2FE6ADBDB5";
    attribute INIT_39 of inst : label is "0BA700BA1EDAA00401955595400A000065555904006AA000410000405A900400";
    attribute INIT_3A of inst : label is "2AFA7ACDA7AB8EFBEBAFA7E8EF23A1E8A6E9E27ED27C702554D14D995508593D";
    attribute INIT_3B of inst : label is "E2F32AAA5705C16EEBAEA7B1FCFEEB7BF0906B3ADDF2ABB7AAEB9EBF2ABAA72F";
    attribute INIT_3C of inst : label is "B92EB0FF67BE7FEB79FBBFA5A7AFB56FB89B9AE8A4AA6ADAB6ABECA94ADAB5AA";
    attribute INIT_3D of inst : label is "D6EA9F9E1DBB2BE1F997F997EAAE197F865FEE4A47E43A0E80EECEDC2B783A6A";
    attribute INIT_3E of inst : label is "1B41D249FA54E292031C33DA6EBFE67EF5ABBFD6FBC6ECAB69FA9FA9CBCAA6BF";
    attribute INIT_3F of inst : label is "901E8AA8E3B8EB9DC89A0BA2496BC93ABEEBB3D6EA7AABF4FFE493BDBFFAF7E4";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
