-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu3 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu3 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "9659D95141A5949DCE826515C425FCF6DAE4B5143C2E5C6A742227D6D60909F4";
    attribute INIT_01 of inst : label is "0D89516965CC2CD7DC9B9A7266535F726E69C9996DA3D893A628D104676545C6";
    attribute INIT_02 of inst : label is "25C5895A925C579A8D7EC083892790D77987690463CC613970A76525467A59FB";
    attribute INIT_03 of inst : label is "88ADE34A8DA424E4A5DE64D27DAE4A55C824B623409F285CC9C97158D8D497BA";
    attribute INIT_04 of inst : label is "1F418481F416960630A0B1E73DB5B9AD69C8DB5388B969289D28289D88D453C8";
    attribute INIT_05 of inst : label is "24548950C619DB18E7E612C85444110961A07D061A07D058481F418481F41848";
    attribute INIT_06 of inst : label is "7F3D65470E7EC5C70676EB373ACD0EB353ACD8EB370257520C9552208494D494";
    attribute INIT_07 of inst : label is "649714252249714AE24E95188D821C52352841C8DA596BD0A35E8DC0A6BB6A0C";
    attribute INIT_08 of inst : label is "DB5B587368B96922263635115C9525266241625A248DC975625A248DC971625A";
    attribute INIT_09 of inst : label is "2523715A95BA23425D56A56E88D09715A958A25C56A5EE89716DE5AE24ED796B";
    attribute INIT_0A of inst : label is "18D04585949E415894854585865A208D66525204141519489C94890505865227";
    attribute INIT_0B of inst : label is "725496888DC58978925C5095B925C56363521A2BB893A545A59473D9A3579097";
    attribute INIT_0C of inst : label is "625C5AA5279F725C5FB893AE8D0001C2F90A35A78898D8D44572549688890545";
    attribute INIT_0D of inst : label is "D8D40585949E572549E417151CEFD654E2725279E625D58949E7989715252791";
    attribute INIT_0E of inst : label is "CD8D8D69A22457254968889050E24E4F6544089CF69672590333DEE7D2FF2E58";
    attribute INIT_0F of inst : label is "2370D89C8DCD8D8D692E245725494A889050E24E95182273DA5906760452743D";
    attribute INIT_10 of inst : label is "88905C96A9250545625494B88DC5CE24E3709486768665117182C8849E67C435";
    attribute INIT_11 of inst : label is "8D86495161A595B5279D84208D6545A59473163635A4A23788A212E45425494B";
    attribute INIT_12 of inst : label is "8D69288DE22C57256208D26C94810545525497888905084D8E24ECD49E747420";
    attribute INIT_13 of inst : label is "87893893A3963635A5A8E274A25A249415154952526237142126CE24ECB9CD8D";
    attribute INIT_14 of inst : label is "7252208DE6C94810508498E24ECD49E7710B3E798D8D69A62457254978889058";
    attribute INIT_15 of inst : label is "2227341F7D253DB6B964E7B21BB9D7412CFFCB98F089422E73E598D8D692E2C5";
    attribute INIT_16 of inst : label is "415256E48DC9755256E48DC9715256249717297BA25C5B49CB893B5272F6D64F";
    attribute INIT_17 of inst : label is "021279A5917102021A592796C509418D051509525E4162521545050652272522";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000008C1C32076F2492FF27795102";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "CB08208208208420821082111082000000000002012301231032230202303210";
    attribute INIT_21 of inst : label is "E772549D5756F96E6A4B78D8DCF86F96EE92F0948D6309CE26584A4941425D74";
    attribute INIT_22 of inst : label is "35C9ED9DEE6372353FFF89FFCB9DEE60B2C124205EF7BAD0522629D89A955457";
    attribute INIT_23 of inst : label is "681D74DE0F0E0F8D2605D5105397FF8FFC9DE7654B73E232773B241C906E6305";
    attribute INIT_24 of inst : label is "D756D35B9ED9D80C0A4589C18985C5C40C008C8884819466919297698A4D4155";
    attribute INIT_25 of inst : label is "1DD5DD1D2AA22AABBB7F0169480000203211194628924891960820B82B5B589A";
    attribute INIT_26 of inst : label is "F6445C65EE8D52557F412F267797F5727440CCCC048C4C40CCCC080888809559";
    attribute INIT_27 of inst : label is "5059BD2357551555554D52F6F4235755055555495CBD690F95117197A3545FC6";
    attribute INIT_28 of inst : label is "C9733346535D04BFC8093929190929059F0D1BA9B257377E154576341548DC8D";
    attribute INIT_29 of inst : label is "A5D84992CE4D24A7D6502517499072B414AD4253B98D755E5233789392919290";
    attribute INIT_2A of inst : label is "AD826DEA5DFFB9297DBB6E054517E7E9FA510509755E4D21092C18BDF48957B9";
    attribute INIT_2B of inst : label is "3753E30151D26576D2F54BE272515571979B7E6942539349A5DE7072B61264B1";
    attribute INIT_2C of inst : label is "24258D77907327B7885549E696509B49CD55543EE11CDC509C111055C63CFED7";
    attribute INIT_2D of inst : label is "030FCCFCEFCDCCCDFDDCDEFC47F54BB614899D424254CDE21567279A59425154";
    attribute INIT_2E of inst : label is "5B716704C31FB38017400CC5CC08DD00331731207400CC0CC089F00321730210";
    attribute INIT_2F of inst : label is "0C300D316DB232CB0FBC05116692EC100813F30C58E01E00C20030C33303FA43";
    attribute INIT_30 of inst : label is "907559249E5A43259D855E6907564949D67676D26189DDCC004C704101E18200";
    attribute INIT_31 of inst : label is "D57195E6907545279690D98B16189D693DA7965B16149D6D37FFFFDE79761C66";
    attribute INIT_32 of inst : label is "9D09D69C77FFFFD279941D5E69279CF41C679082696109D693DE79A584275299";
    attribute INIT_33 of inst : label is "BB6652642779925C6549E79A5A41507571279C8527537FFFD9555690C9F961E9";
    attribute INIT_34 of inst : label is "587195D79A42DC71A9C2A41D5D49E43D072B9C4A655675365842743CCAE536FD";
    attribute INIT_35 of inst : label is "7649C899F06A9FE69C655472A79A5D16E49C999F0629F2790755472649E58427";
    attribute INIT_36 of inst : label is "4275A710A984D77FFFDDA67195E79A7D072B94B71CAA41D5D49E70A96109D6D1";
    attribute INIT_37 of inst : label is "07549E79A4D77FFFE9943655CD5365A43E587E427535DFFDD265A4365E586A67";
    attribute INIT_38 of inst : label is "9719988A596109D511641C069C19C1CA9C1C6579A59271967040E9CD9C1C29D1";
    attribute INIT_39 of inst : label is "00F3FCDCDCFCFCDC10DC10DC10DC10DC0FC303010303030102F4D77FFE75365D";
    attribute INIT_3A of inst : label is "0F1C2D3E0F004073C3C340B400000003CCC0C0C3E3E1D1D00C0C0C0C0B000000";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF33D5D1011912C3C7434073E2D1C";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "F5E6B5D7807D746B8BAF7E79201F42ADB37DD31018F7E2F3E7317EB9BBA7275C";
    attribute INIT_01 of inst : label is "3B65D79F5FB8EC9E366479F997C278D951E7E55F9BF2B0B93C84B0009AD75EC1";
    attribute INIT_02 of inst : label is "A70328EF6A7139FF49EA91EB6F7C73B5EF65EF89CBADC3A7969F7F975CD7D7AA";
    attribute INIT_03 of inst : label is "4C5BB9C24B2C9C5C5D717D77C713C1CD44B02D92FAFE0A726FE9C4E4B4B88DD4";
    attribute INIT_04 of inst : label is "0BE86C4CBE893D20A9DB577FAB6CDFF4C804B12103DF93F2EBBA7EEB84B9F119";
    attribute INIT_05 of inst : label is "8EA846B2DC1729701C6A2BA4C70002079B112F81B102F826C4CBE86C44BE86C4";
    attribute INIT_06 of inst : label is "87FFA79CB1C6B79CB5CA082D8E3B228AE861B2082E98EAA1A23AA11A623AA86B";
    attribute INIT_07 of inst : label is "5A9C0CA3BDA9C4DC13C25D76CB4FEC1B2DAF80CCB7D74AB612D8CB0011331100";
    attribute INIT_08 of inst : label is "B6CD362142DF93D3192D2E81B68DA79BD210FA37984BE9C8DA37984BE9C8FA37";
    attribute INIT_09 of inst : label is "A7D20CDAACC612CA7236AB3184B29C8DAACC6A7036AB35A9C4EF7DC13C2ADF4A";
    attribute INIT_0A of inst : label is "74B64B60AFF7C0529E4C730BA2B756CB755A7921CF2C8ADE5A9E4843CBE2BB96";
    attribute INIT_0B of inst : label is "CA369FF74833A8DD6A703E8EE6A71392F2EA375604F0975E7D702AB512E44079";
    attribute INIT_0C of inst : label is "3A7036A3FDF43A713404F0AC4B0006185F6B2E4C5C64B4BA06DA369EF6484306";
    attribute INIT_0D of inst : label is "B4BA8B688FF7DBA7BF7C0A3B7657063253FA3FDF03A72368FF7C0E9C8FA3FDF0";
    attribute INIT_0E of inst : label is "A24B4B9357106FA369EF64843C13C2AAD75D8F342DF5EAAAADD1693941FF17E4";
    attribute INIT_0F of inst : label is "B2EB2A7CCBA24B4B93DF106FA369EE64843C13C25D7A7CD0B7D7C7CAA9D1ADAB";
    attribute INIT_10 of inst : label is "6484368EF6A74306FA369FF74833013C2ACA74A7CA01BE75C76BA2F9F1CD00ED";
    attribute INIT_11 of inst : label is "CBABF5D7807D79A77C7A00E0CB975E7D700B092D2E4FCB2C6C5237506CA369EF";
    attribute INIT_12 of inst : label is "4B93F2CB1B106DA3BD6CBBD29E487306FA369DC6484388E0813C2E9DF1E86CE6";
    attribute INIT_13 of inst : label is "8CD504F08A392D2E4F4E8BAC4A379A9D0C1BA8DA7B9D20CD2331413C2AA3A24B";
    attribute INIT_14 of inst : label is "FA3B96CB7929E487348D0C13C2A9DF1E803A87EE4B4B9313106FA369DF648438";
    attribute INIT_15 of inst : label is "8BBE8A78E0BFAB6CDFB67ED39D5F4EB41CDFC5F053EF2317E87EE4B4B93D3106";
    attribute INIT_16 of inst : label is "10DAB3184BE9C8FAB3184BE9C8DAB31A9C0E2ACD6A713BEF904F0ABBEAADB346";
    attribute INIT_17 of inst : label is "E3EFE77D75C74BABEBE77C7B8007A74B692EAACFD7C08A793273CBE2B796A792";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000001102549B313B01FF1995D783";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "3B00000000000000000000000000004010040120321003211330211003220321";
    attribute INIT_21 of inst : label is "92F07A4B377400C033C43CB4BA61C00C04F130764B4407413C8801F4F0C0F33F";
    attribute INIT_22 of inst : label is "0044DDF453F6EB6C91545FFFC4F4D3F8F14016301311BFE0213C2CB00CF3921F";
    attribute INIT_23 of inst : label is "3001CC456EAD46DB7C1733601105547FFC74DF848749D917CD377C017001C08B";
    attribute INIT_24 of inst : label is "F2F2F2B67AFA727A76723EB2763A727A7E767A727A720C5CF31075CF87B38403";
    attribute INIT_25 of inst : label is "004C084CC88C04C8448C814848203211000020C3C86D04F07904003E7CFCFF32";
    attribute INIT_26 of inst : label is "1ECF39E731CBB30DF380123F2DC301E32C8CC048048C4808C4C4084C8400CCCC";
    attribute INIT_27 of inst : label is "7716CB32CCBB21CCDEC47B2D2D32CCBB11CCDECC724B8F44FB3CE79CF2EC8E23";
    attribute INIT_28 of inst : label is "4F66664656AE707FC7170707070717A439393646658D0CC0825C752C07A4BACB";
    attribute INIT_29 of inst : label is "8E34CC7345E7FC5E73D85D77CC7009EC0CFB81D37F4B1DBDD061F7F070707178";
    attribute INIT_2A of inst : label is "CB4DC7DFC7577F07A7C9F2B74579BC6F1FD7DE279DBDD75E0750767B484F1F7F";
    attribute INIT_2B of inst : label is "AA83A9806DF3DC7841DE871DDFE307B7DE38F9EF81E075FF4D38F01B2D331CD7";
    attribute INIT_2C of inst : label is "1C1E4B1EF0C93D9F71C7973C73E079CF8DE31E2A98AAA6B63E880037291A6AA0";
    attribute INIT_2D of inst : label is "0895645645467467546464658C01C4F9084FCB81C5EE47DC71CF5CF1CF81D178";
    attribute INIT_2E of inst : label is "3B706704C3073182B3C00C43C4068F00310F001B3C00C40C406CF00310F101B0";
    attribute INIT_2F of inst : label is "0CB2C002A08331C10C30A083F0C3CC92CF3BE18EF861BF40C20033C23105F983";
    attribute INIT_30 of inst : label is "F5C7977D73E3D1BE4B9E71CF5C71CFE4B92D2C7BD70CBCC4080C308000208308";
    attribute INIT_31 of inst : label is "B9D75E5DF5C7885CF8F46FA6F178CB8F079C7BE6F178CBB79FBBBB75FF9E709D";
    attribute INIT_32 of inst : label is "4BCCB8F05FBBB97DDF5D71E9EF5CF21D709CF22BDF974CB8F075C77E5D32E474";
    attribute INIT_33 of inst : label is "C9FA81FCFDC7F275D7B7BD77E3D275C7B05CFA5D32E9FBBBAF9E78F46FC79787";
    attribute INIT_34 of inst : label is "E9D75EF177C975C25FC3BD71EE173C875C34FE2FBE7B2D1BE5D32CFC45D6DF27";
    attribute INIT_35 of inst : label is "A6A3C4F3E0203EDFF5D792A1BD77E77A6A3C7F3E0243EDEF5C792A1BD73E5D32";
    attribute INIT_36 of inst : label is "F32E3C98EF9E75FBBBA7DBD75EF177C75C04FE5D7017D71EF173F0EF974CBA77";
    attribute INIT_37 of inst : label is "5C7973E7BE75FBBBBFDD97E76DD1BE3D1FE5FDE32E9D7FF679BE3D17C1E5E1D2";
    attribute INIT_38 of inst : label is "9C06F209EF974CBB7DCC0FB23FC3C0B83C05D7977F7FE79CF03B63C03C0B03C0";
    attribute INIT_39 of inst : label is "00F1141414040414581458145814581401404C014D0C0C0D00CA75FFDBE797E7";
    attribute INIT_3A of inst : label is "31323232020073503030703400000003C5425251414252502525141403000000";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF11DDD1015550C3C570406323232";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "924C134D412496C1733F34D3B8370330C1014815A7334BF3403A7CC0C10D0F3E";
    attribute INIT_01 of inst : label is "B6134D451532EA100780131E0378401E004C780D0C14C0CA34881000304D35C4";
    attribute INIT_02 of inst : label is "84AB70000849B00130130CC9AF249B634D134D3C8B308D85CA14364D35A2494C";
    attribute INIT_03 of inst : label is "500C136B01103D3C3CF134F34F1343EECD3200404CD8ACD68D6126C838130011";
    attribute INIT_04 of inst : label is "820D004423D0011048C88D36CC3040120120105A04CD00424141424120135D9C";
    attribute INIT_05 of inst : label is "D968499F08C59C231673530019B0000D0013080401308C400482010048231004";
    attribute INIT_06 of inst : label is "2AEB0F3CD1678F3CD16718584206508194206908195DAA626F65A1269F6A989A";
    attribute INIT_07 of inst : label is "4212AEC0002126C4226334D1813FDC5605CF4128124904C22040410002112000";
    attribute INIT_08 of inst : label is "C314804A06CD0018020E047A730084200062DC000203212EFC000203212ACC00";
    attribute INIT_09 of inst : label is "84006ECD300080D84BB34C00203612ACD301084AB34C002126C434C226320D04";
    attribute INIT_0A of inst : label is "D83197313003C04610019B97B0C00243001840066E5DC3000210018B97B0C000";
    attribute INIT_0B of inst : label is "EC02100081BBF001084AB30000849B20604880020898CD351450ACC3204EE0D0";
    attribute INIT_0C of inst : label is "084AB34000D00849B00898C4814103088D22040060083811E9CC021000818BE9";
    attribute INIT_0D of inst : label is "381197340003C484403407B72213DAB2237C000D0084BB7000340212AEC000D4";
    attribute INIT_0E of inst : label is "00818300140E9CC021000818B62263F30D34CF6A989240C80080A9946140E348";
    attribute INIT_0F of inst : label is "507F9CC24100818300180E9CC021000818B6226334DF3DAA62493367134A06CC";
    attribute INIT_10 of inst : label is "0818BF0000849BE9CC02100081BB62263304C323676234D34D3307F4515A0ADB";
    attribute INIT_11 of inst : label is "4173734D41249040249906EE410D3524904712060C0209046018800E9EC02100";
    attribute INIT_12 of inst : label is "8300824118CA9DC00024300610819BE9FC021010818B620022263B0092669AE5";
    attribute INIT_13 of inst : label is "20028898CC42060C00720B041C0002126FA7B008400206EC8800E22630440081";
    attribute INIT_14 of inst : label is "CC00024300610819BE200A226330092641B800048183001C0E9CC021000818BA";
    attribute INIT_15 of inst : label is "1B3400D10A34CC3140110048CC8D224E140038DE8CCD67E3400048183001C0A9";
    attribute INIT_16 of inst : label is "62CCC00203212EDCC00203212AFCC04212AC13000849B10D00898C834130C528";
    attribute INIT_17 of inst : label is "33D24914534DBFB3D2491453220D0D83165D332023C05840059B97B0C0008400";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFE010C10C300300000000003834A140E3234D33";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "17410410E104010E380438000438EE3B8EE3B844777776666556555554444777";
    attribute INIT_21 of inst : label is "B048D2C19891051033CEC0101603D05108F380D641900D2235A403E262F85174";
    attribute INIT_22 of inst : label is "06D028DC23704B0570008D4038DC235AC002133CAB843F1462250C140CFB842C";
    attribute INIT_23 of inst : label is "4023E7C22C1C2CC1348F980AAFE000B803B42C558AA73CA3640A3500FC83D095";
    attribute INIT_24 of inst : label is "E5A1EDE925E121A5A96DA1A1EDA9292521A1A9A5ADA8500CF500F3CF23C94189";
    attribute INIT_25 of inst : label is "048C4804C4C4080C840CC0484A110000000005038CD88450D3E03CDDA9E1E9A9";
    attribute INIT_26 of inst : label is "353CF3CF88C3302E485218160542AA5A04CCC000444488CCC00488CC048CC048";
    attribute INIT_27 of inst : label is "B6800130E5C50666E54D900404B0E5C50666E5419A011428D0F3CF3E30DC9243";
    attribute INIT_28 of inst : label is "9F666664762168503B0D0D0D0D0D0FD620B1C647772D6EE84A55430D8F2C36C3";
    attribute INIT_29 of inst : label is "7DF5003287DF3C3DF3E43CF604700B0CC6C3034B8FC33D42D0C348F0D0D0D0F6";
    attribute INIT_2A of inst : label is "8331DF23DF008F0F0FE3F85F2D033ECFB3D07C0F3D42CD3C1F71F2C3E457A78F";
    attribute INIT_2B of inst : label is "6A4F0AC24D811C85E14C0014C7C12B0F3CF3C2CB03C1F7CF7DF9A08A0D404CA2";
    attribute INIT_2C of inst : label is "3C34C33CF34A343CB7DF575DB6C0F3DF23CB6ED30BD30D7329BC10BBD7E09337";
    attribute INIT_2D of inst : label is "0547665446775547776647543956420558898103C3468D2DF7DA5D76DB03C9F0";
    attribute INIT_2E of inst : label is "224034000003000033C000020014CF22C00800173C8B0000005CF22C00800150";
    attribute INIT_2F of inst : label is "A04111440104C000308210400000C0830C31C00C90003F5E0000C108C000FD78";
    attribute INIT_30 of inst : label is "D34D555492450A348134D65934D65968120704D75C681C0003208212480208CC";
    attribute INIT_31 of inst : label is "134D3524934D412491428D9499C281140D24134499C2810D373330D44D34D305";
    attribute INIT_32 of inst : label is "C1281142373330D04D34D34041249534D304D6734D1C281140D2413470A040DC";
    attribute INIT_33 of inst : label is "E37521153340D0D34D4514924508D34D79249D70A04373330D34D1428D0D1C0D";
    attribute INIT_34 of inst : label is "434D34F09254D34C0D3734D34F09254D34D0D27F34D204A3470A04FF00F0378D";
    attribute INIT_35 of inst : label is "D3268556A05F6A14534D02C004924D2D3268456A05F6A14534D02C00492470A0";
    attribute INIT_36 of inst : label is "4A04508DCD34D373330DC34D35F4924D34C0D534D3034D35F4925DCD1C2810D2";
    attribute INIT_37 of inst : label is "34D0924104D373330D35A34D934A3450A347334A0434D558D13450A343470370";
    attribute INIT_38 of inst : label is "34C4DD234D1C2810D348289B6816829368934D0924104D34A089B68D68297689";
    attribute INIT_39 of inst : label is "00F0848484848484848484848484848488484448444444444400D355634D234D";
    attribute INIT_3A of inst : label is "11111111212211121212110000000003C0101010101010120101010110000000";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF04000484444403C112221111111";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "71F8F1C7081C704F0B071C3C700CF01CF00C03602031F0F1CB771C7CF003031D";
    attribute INIT_01 of inst : label is "5741C7071CCD400C37CCB3DF31C030DF32CF7CC7CF0C77C21D34F000F3C71CE0";
    attribute INIT_02 of inst : label is "035301C000353C3002CCC0C0C71C7571C701C709C1D5C00B502D1C071DE1C733";
    attribute INIT_03 of inst : label is "130F01DCCF7C0D0C0C731C71C731C0FF6E047D23D0B370308740D4FCFCF01C00";
    attribute INIT_04 of inst : label is "83CC0C383FCC30E100C0C31D073C0300DC04F7027CC7C3404F40404F04F0C050";
    attribute INIT_05 of inst : label is "1D0001425C0B51702D4F0DC004000303C30F0F0030F0FC30C3C3C00C383F00C3";
    attribute INIT_06 of inst : label is "C451C71D72D4C71D72D4619C18670619C18670619C01C700507400050071C014";
    attribute INIT_07 of inst : label is "000D4D070000D4D732D01C708F074E033C2D0804F1C76C75D3DB4F0030000300";
    attribute INIT_08 of inst : label is "73C035026CC7C304CF3F3C30301C03000018C070004F00D4C070004F00D4D070";
    attribute INIT_09 of inst : label is "03001CD70C0013C03535C30004F00D4D70C0003535C30000D4C31D732D02C76C";
    attribute INIT_0A of inst : label is "3CF0C30F0D31C0F00C0043C30C30004F00C03001CF0D30C0300C0063C34C300C";
    attribute INIT_0B of inst : label is "C0700C00007301C00035341C000353F3F3C07004CCB4071C1C703074D3F1C03C";
    attribute INIT_0C of inst : label is "003537C74C70003534CCB41B4F4105D7875D3F0C133CFCF0C0C0700C000063C0";
    attribute INIT_0D of inst : label is "FCF0C30F1D31FC03D31C0F037037C53431C074C700035341D31C000D4D074C70";
    attribute INIT_0E of inst : label is "7FCFCFC300CC0C0700C000063032D001C71D1D79DC71DD1D9DD93D11004071FC";
    attribute INIT_0F of inst : label is "33D251B04F7FCFCFC3048C0C0700C000063032D01C7075E771C742D400C13D07";
    attribute INIT_10 of inst : label is "0006301C000373C0D0700C000073432D06C1B002D4031C31C7037FD071DE315D";
    attribute INIT_11 of inst : label is "CF02D1C7001C76CB1C7C01404FC71C1C70030F3F3F0C013C0300700C0C0700C0";
    attribute INIT_12 of inst : label is "CFC3004F00CC0C070004F0000C0073C0C0700C00006341C0432D042C71F1DD40";
    attribute INIT_13 of inst : label is "1C000CB411FF3F3F0C13C13E0070000DCF0301C0300001CD0700032D07DF7FCF";
    attribute INIT_14 of inst : label is "C070004F0000C007301C0032D042C71F0051F0C3CFCFC3048C0C0700C0000630";
    attribute INIT_15 of inst : label is "F31DFC32C81C073C03000C000CC70F1006101C7090C74371DF0C3CFCFC3048C0";
    attribute INIT_16 of inst : label is "18D030004F00D4D030004F00D4D030000D4DF0C0003530C77CCB40B1DF1CF009";
    attribute INIT_17 of inst : label is "0741C71C71C70F0341C71C7FD003C3CF0F0F00F4F1C0C0300343C30C300C0300";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFF01001000000000000000D919100407CE1C70F";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "1B00000000000000000000000514501405014066555555555555555555555444";
    attribute INIT_21 of inst : label is "E3C0304FFFFD36D331E07CF8F070D36D387030304FD303031D0000D0D0C06174";
    attribute INIT_22 of inst : label is "034E307631E3C13C1800C7403C7631C3DBB070783116FDC4001D34F4CC7FF43F";
    attribute INIT_23 of inst : label is "6F00CD63070C078F1F033D40357800D403D6371C01C13421CD8C1E803800D383";
    attribute INIT_24 of inst : label is "559551511151119D9D1D1D9D59191919D999151511136F2C76C031C7034300FF";
    attribute INIT_25 of inst : label is "444488CCC00488CC0488C04848000000000836F3400400703F0F0821911D1555";
    attribute INIT_26 of inst : label is "1C1C71C711CF303FF310031F3F420FD13C0004444444444448888888CCCCC000";
    attribute INIT_27 of inst : label is "F4038FD3FDF303FFFCC0FD3E3C13FDF303FFFCC0F04FDB087C71C71C73CC0F33";
    attribute INIT_28 of inst : label is "8765555545FC50101D03030303030304DC1DB66544FF0CC03FD0FE3C0304F04F";
    attribute INIT_29 of inst : label is "1C74C07040C71E0C71C30C77C072013CC04FC0C0C7CF1DF35371CC7030303030";
    attribute INIT_2A of inst : label is "CF02C731C700C783C741D00301FD1C4711DF0FC31DF347F7034C304F4007FCC7";
    attribute INIT_2B of inst : label is "3300C240F5F01FF180630132E1C03FC71C71F1C7C0F031C71C7DE0013D301C17";
    attribute INIT_2C of inst : label is "0C0FCF1C71C21D1CD1C7071C71F031C700FFFF0CC24CCC307824003FC30F8CDF";
    attribute INIT_2D of inst : label is "044777777666666555555444EC0FC071C007CFC0C0FC873471DE1C71C7C0C03C";
    attribute INIT_2E of inst : label is "2240340104020C0033C0B3023000CF11CC08C0033C473003020CF11CC08C0840";
    attribute INIT_2F of inst : label is "A082030C030CCC0030C20104010440C00010CC0CF3003F9D00000200CC00FD74";
    attribute INIT_30 of inst : label is "71C7071C71F6C21F8F1C71C71C71C704FF3F3C71DB04FC3003104100000000C0";
    attribute INIT_31 of inst : label is "F0C71C1C71C7001C7DB0870F41B04FDBC72CB1FF41B04FC71CCCCC72C71C302C";
    attribute INIT_32 of inst : label is "CF04FDB01CCCCC72C70C71C1C71C701C302C7002C7DB04FDBC72CB1F6C13F03C";
    attribute INIT_33 of inst : label is "41D1001F31CC7C31C7071C71F6C031C73C1C706C13F1CCCCC70C3DB08703DB03";
    attribute INIT_34 of inst : label is "F0C71CF071C070C0C7031C71CF071C070C0C70031C3E3C21F6C13C7F00F31D07";
    attribute INIT_35 of inst : label is "53078077B01F7B1C71C700701C71C775F078077B01B7B1C71C700701C71F6C13";
    attribute INIT_36 of inst : label is "C13F6C01C70C71CCCCC7F1C71CF071C70C0C701C3031C71CF071C0C7DB04FC77";
    attribute INIT_37 of inst : label is "1C7071C71C71CCCCC70C21C3C0C21F6C21F6F0C13F1C7008731F6C21C0F6C0F3";
    attribute INIT_38 of inst : label is "0C0C7C02C7DB04FC71DC081778C780D77841C7071C71C71DE0013780780D3780";
    attribute INIT_39 of inst : label is "00F004141404041414141414141414148040404140404041480C71C021C3E1C7";
    attribute INIT_3A of inst : label is "01010101012090901010920000000003C0909090909090920909090920000000";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF02111182222803C090505010101";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
