library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_PROG_ROM_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_PROG_ROM_2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"A5",X"17",X"49",X"FF",X"A8",X"A5",X"18",X"49",X"FF",X"AA",X"C8",X"D0",X"01",X"E8",X"98",X"18",
		X"65",X"1B",X"A8",X"8A",X"A2",X"00",X"65",X"1C",X"10",X"05",X"98",X"49",X"FF",X"A8",X"CA",X"86",
		X"40",X"60",X"20",X"F9",X"6F",X"98",X"A4",X"3D",X"20",X"C0",X"70",X"A5",X"1D",X"38",X"E5",X"15",
		X"A4",X"77",X"20",X"EF",X"70",X"86",X"37",X"A4",X"76",X"20",X"F1",X"70",X"18",X"65",X"37",X"85",
		X"37",X"24",X"40",X"30",X"0E",X"18",X"65",X"17",X"85",X"48",X"A5",X"18",X"69",X"00",X"85",X"49",
		X"4C",X"60",X"70",X"38",X"A5",X"17",X"E5",X"37",X"85",X"48",X"A5",X"18",X"E9",X"00",X"85",X"49",
		X"A6",X"1F",X"A5",X"20",X"20",X"9B",X"70",X"10",X"04",X"A2",X"8F",X"86",X"5D",X"60",X"20",X"F9",
		X"6F",X"A5",X"3D",X"20",X"C0",X"70",X"A5",X"17",X"38",X"E5",X"1F",X"A4",X"77",X"20",X"EF",X"70",
		X"86",X"37",X"A4",X"76",X"20",X"F1",X"70",X"18",X"65",X"37",X"85",X"37",X"18",X"65",X"15",X"85",
		X"48",X"A5",X"16",X"69",X"00",X"85",X"49",X"A6",X"1D",X"A5",X"1E",X"85",X"4B",X"A9",X"80",X"24",
		X"49",X"10",X"14",X"A5",X"48",X"49",X"FF",X"85",X"48",X"A5",X"49",X"49",X"FF",X"85",X"49",X"E6",
		X"48",X"D0",X"02",X"E6",X"49",X"A9",X"00",X"85",X"4C",X"A0",X"00",X"84",X"4D",X"4C",X"02",X"6D",
		X"84",X"75",X"20",X"D1",X"70",X"86",X"77",X"A2",X"00",X"86",X"78",X"20",X"D5",X"70",X"86",X"76",
		X"60",X"85",X"78",X"A9",X"00",X"A0",X"07",X"26",X"78",X"2A",X"B0",X"0E",X"C5",X"75",X"90",X"02",
		X"E5",X"75",X"88",X"10",X"F2",X"26",X"78",X"A6",X"78",X"60",X"E5",X"75",X"38",X"B0",X"F3",X"85",
		X"43",X"84",X"42",X"A5",X"43",X"48",X"49",X"FF",X"85",X"43",X"A9",X"00",X"85",X"44",X"85",X"45",
		X"A2",X"08",X"06",X"43",X"B0",X"06",X"65",X"42",X"90",X"02",X"E6",X"45",X"CA",X"D0",X"07",X"AA",
		X"68",X"85",X"43",X"A5",X"45",X"60",X"0A",X"26",X"45",X"90",X"E7",X"55",X"A9",X"00",X"85",X"55",
		X"85",X"57",X"A9",X"0F",X"24",X"4E",X"50",X"02",X"A9",X"03",X"85",X"37",X"A5",X"08",X"24",X"5A",
		X"10",X"0D",X"C9",X"20",X"B0",X"1A",X"20",X"2C",X"73",X"B0",X"15",X"C6",X"4F",X"90",X"0B",X"C9",
		X"E0",X"90",X"0D",X"20",X"1B",X"73",X"90",X"08",X"E6",X"4F",X"A5",X"4F",X"25",X"37",X"85",X"4F",
		X"24",X"4E",X"50",X"03",X"4C",X"3E",X"72",X"A5",X"0A",X"24",X"5C",X"10",X"0A",X"C9",X"40",X"B0",
		X"03",X"20",X"54",X"73",X"4C",X"03",X"72",X"C9",X"A5",X"90",X"F9",X"20",X"FE",X"72",X"C9",X"02",
		X"90",X"06",X"D0",X"0A",X"E0",X"08",X"B0",X"06",X"20",X"3D",X"73",X"4C",X"03",X"72",X"24",X"5D",
		X"10",X"03",X"4C",X"39",X"72",X"A5",X"0F",X"18",X"65",X"51",X"85",X"51",X"A5",X"10",X"29",X"03",
		X"65",X"4F",X"29",X"0F",X"AA",X"4A",X"66",X"51",X"4A",X"66",X"51",X"18",X"69",X"02",X"29",X"03",
		X"85",X"4F",X"8A",X"29",X"0C",X"48",X"0A",X"0A",X"AA",X"BD",X"E2",X"51",X"38",X"E5",X"53",X"85",
		X"48",X"BD",X"E3",X"51",X"E5",X"54",X"85",X"49",X"A9",X"80",X"85",X"4C",X"A0",X"00",X"A6",X"0D",
		X"A5",X"0E",X"29",X"0F",X"20",X"FE",X"6C",X"4A",X"66",X"4A",X"4A",X"66",X"4A",X"85",X"4B",X"68",
		X"AA",X"BD",X"BC",X"4B",X"85",X"48",X"BD",X"BD",X"4B",X"85",X"49",X"A9",X"00",X"85",X"50",X"85",
		X"52",X"85",X"53",X"85",X"54",X"85",X"09",X"85",X"07",X"85",X"4C",X"20",X"04",X"6D",X"84",X"0A",
		X"4A",X"66",X"0A",X"66",X"09",X"4A",X"66",X"0A",X"66",X"09",X"A9",X"80",X"85",X"08",X"A9",X"40",
		X"85",X"4E",X"60",X"20",X"FE",X"72",X"09",X"00",X"D0",X"2B",X"E0",X"02",X"B0",X"27",X"C0",X"02",
		X"B0",X"23",X"A5",X"02",X"38",X"E9",X"07",X"C9",X"03",X"B0",X"1E",X"A5",X"61",X"A2",X"80",X"C9",
		X"04",X"90",X"06",X"C9",X"08",X"B0",X"12",X"A2",X"C0",X"A5",X"5F",X"C9",X"04",X"B0",X"0A",X"8A",
		X"05",X"5D",X"85",X"5D",X"60",X"24",X"5D",X"10",X"04",X"A9",X"8F",X"85",X"5D",X"60",X"A5",X"0A",
		X"24",X"5C",X"30",X"1A",X"C9",X"A5",X"90",X"2A",X"20",X"3D",X"73",X"F0",X"10",X"C9",X"02",X"90",
		X"0C",X"20",X"2D",X"65",X"20",X"96",X"6B",X"A2",X"FF",X"9A",X"4C",X"40",X"60",X"60",X"A5",X"53",
		X"05",X"54",X"F0",X"0E",X"20",X"54",X"73",X"B0",X"F4",X"A9",X"00",X"85",X"52",X"85",X"53",X"85",
		X"54",X"60",X"20",X"FE",X"72",X"A8",X"D0",X"F9",X"E0",X"60",X"B0",X"F5",X"A5",X"0F",X"18",X"65",
		X"51",X"85",X"51",X"A5",X"10",X"65",X"4F",X"29",X"03",X"AA",X"06",X"51",X"2A",X"06",X"51",X"2A",
		X"48",X"38",X"E9",X"02",X"29",X"0F",X"85",X"4F",X"8A",X"0A",X"0A",X"AA",X"BD",X"BC",X"4B",X"85",
		X"48",X"BD",X"BD",X"4B",X"85",X"49",X"A9",X"80",X"85",X"4C",X"A5",X"0E",X"A6",X"0D",X"A0",X"00",
		X"20",X"FE",X"6C",X"06",X"4A",X"2A",X"06",X"4A",X"2A",X"85",X"4B",X"A9",X"A3",X"A2",X"78",X"85",
		X"49",X"86",X"48",X"20",X"04",X"6D",X"A9",X"18",X"85",X"48",X"A9",X"A1",X"85",X"49",X"A9",X"00",
		X"85",X"4C",X"85",X"4E",X"85",X"07",X"85",X"09",X"85",X"50",X"85",X"52",X"20",X"04",X"6D",X"68",
		X"29",X"0C",X"0A",X"AA",X"BD",X"22",X"52",X"85",X"48",X"BD",X"23",X"52",X"85",X"49",X"20",X"04",
		X"6D",X"85",X"54",X"84",X"53",X"A9",X"80",X"85",X"08",X"A9",X"9E",X"85",X"0A",X"60",X"A0",X"FF",
		X"A5",X"7E",X"A6",X"7D",X"C5",X"80",X"90",X"12",X"D0",X"0C",X"A4",X"7F",X"C4",X"7D",X"B0",X"0A",
		X"A6",X"7F",X"A4",X"7D",X"90",X"04",X"A5",X"80",X"A6",X"7F",X"60",X"20",X"6B",X"73",X"A5",X"50",
		X"18",X"65",X"3D",X"85",X"50",X"A5",X"51",X"65",X"3E",X"85",X"51",X"60",X"20",X"6B",X"73",X"A5",
		X"50",X"38",X"E5",X"3D",X"85",X"50",X"A5",X"51",X"E5",X"3E",X"85",X"51",X"60",X"20",X"8A",X"73",
		X"A5",X"52",X"18",X"65",X"3F",X"85",X"52",X"A5",X"53",X"65",X"40",X"85",X"53",X"A5",X"54",X"69",
		X"00",X"85",X"54",X"60",X"20",X"8A",X"73",X"A5",X"52",X"38",X"E5",X"3F",X"85",X"52",X"A5",X"53",
		X"E5",X"40",X"85",X"53",X"A5",X"54",X"E9",X"00",X"85",X"54",X"60",X"A9",X"80",X"85",X"55",X"A5",
		X"5F",X"85",X"3D",X"A9",X"00",X"85",X"3E",X"A5",X"5E",X"A2",X"02",X"24",X"4E",X"70",X"02",X"A2",
		X"04",X"0A",X"26",X"3D",X"26",X"3E",X"CA",X"D0",X"F8",X"60",X"A9",X"80",X"85",X"57",X"A5",X"61",
		X"85",X"3F",X"A9",X"00",X"85",X"40",X"A5",X"60",X"A2",X"02",X"24",X"4E",X"70",X"02",X"A2",X"04",
		X"0A",X"26",X"3F",X"26",X"40",X"CA",X"D0",X"F8",X"60",X"A9",X"BA",X"85",X"64",X"A9",X"51",X"85",
		X"65",X"A9",X"45",X"85",X"28",X"A9",X"6B",X"85",X"69",X"A9",X"00",X"85",X"27",X"85",X"6A",X"85",
		X"37",X"85",X"38",X"85",X"39",X"A9",X"F0",X"85",X"2B",X"A9",X"44",X"85",X"2C",X"20",X"03",X"75",
		X"A0",X"00",X"B1",X"64",X"AA",X"C8",X"B1",X"64",X"C9",X"A0",X"90",X"12",X"C9",X"D0",X"90",X"25",
		X"F0",X"4F",X"91",X"27",X"88",X"8A",X"49",X"08",X"91",X"27",X"C8",X"C8",X"D0",X"E4",X"38",X"E9",
		X"20",X"91",X"27",X"88",X"8A",X"91",X"27",X"C8",X"C8",X"B1",X"64",X"91",X"27",X"C8",X"B1",X"64",
		X"91",X"27",X"C8",X"D0",X"CD",X"29",X"0F",X"85",X"3A",X"86",X"3B",X"88",X"20",X"F8",X"74",X"C8",
		X"C8",X"98",X"A0",X"00",X"18",X"65",X"64",X"91",X"69",X"E6",X"69",X"A5",X"65",X"69",X"00",X"91",
		X"69",X"E6",X"69",X"A5",X"3B",X"0A",X"85",X"64",X"A5",X"3A",X"2A",X"09",X"40",X"85",X"65",X"D0",
		X"A1",X"88",X"20",X"F8",X"74",X"A0",X"00",X"C6",X"69",X"B1",X"69",X"85",X"65",X"C6",X"69",X"B1",
		X"69",X"85",X"64",X"A6",X"69",X"E0",X"6B",X"D0",X"89",X"E6",X"37",X"A2",X"04",X"E4",X"37",X"D0",
		X"81",X"A9",X"00",X"85",X"37",X"91",X"27",X"C8",X"A9",X"D0",X"91",X"27",X"C8",X"20",X"F8",X"74",
		X"E6",X"39",X"A2",X"04",X"E4",X"39",X"F0",X"03",X"4C",X"CD",X"73",X"A9",X"F0",X"85",X"64",X"A9",
		X"44",X"85",X"65",X"A5",X"38",X"18",X"65",X"2B",X"85",X"2B",X"D0",X"02",X"E6",X"2C",X"A0",X"07",
		X"B1",X"64",X"91",X"2B",X"88",X"10",X"F9",X"A9",X"7E",X"85",X"64",X"A9",X"4E",X"85",X"65",X"A9",
		X"00",X"85",X"27",X"A9",X"47",X"85",X"28",X"A0",X"00",X"A2",X"00",X"B1",X"64",X"E0",X"01",X"D0",
		X"05",X"38",X"E9",X"20",X"D0",X"16",X"E0",X"07",X"D0",X"12",X"29",X"03",X"85",X"37",X"88",X"B1",
		X"64",X"46",X"37",X"6A",X"46",X"37",X"6A",X"91",X"27",X"C8",X"A9",X"04",X"91",X"27",X"E8",X"8A",
		X"29",X"07",X"AA",X"C8",X"C0",X"20",X"90",X"D3",X"A5",X"21",X"F0",X"2B",X"A2",X"05",X"86",X"37",
		X"0A",X"AA",X"CA",X"CA",X"A9",X"40",X"85",X"27",X"A9",X"47",X"85",X"28",X"BD",X"6A",X"5E",X"BC",
		X"69",X"5E",X"20",X"A4",X"7E",X"A6",X"65",X"A4",X"64",X"20",X"F2",X"79",X"A5",X"2C",X"A4",X"2B",
		X"20",X"CD",X"7E",X"C6",X"37",X"10",X"EE",X"60",X"98",X"18",X"65",X"27",X"85",X"27",X"90",X"02",
		X"E6",X"28",X"60",X"A5",X"28",X"4A",X"29",X"0F",X"09",X"C0",X"AA",X"A5",X"27",X"6A",X"A4",X"38",
		X"91",X"2B",X"8A",X"C8",X"91",X"2B",X"C8",X"84",X"38",X"60",X"A8",X"A2",X"03",X"86",X"39",X"A2",
		X"02",X"B5",X"5F",X"B4",X"5E",X"84",X"37",X"A0",X"09",X"86",X"3A",X"AA",X"20",X"C6",X"79",X"48",
		X"8A",X"A6",X"39",X"95",X"A7",X"94",X"A8",X"68",X"95",X"A6",X"A6",X"3A",X"A0",X"02",X"05",X"94",
		X"05",X"93",X"F0",X"07",X"B5",X"5A",X"0A",X"A9",X"00",X"2A",X"A8",X"8A",X"4A",X"AA",X"94",X"9A",
		X"A9",X"00",X"85",X"39",X"A6",X"3A",X"CA",X"CA",X"10",X"C7",X"20",X"FE",X"72",X"86",X"37",X"24",
		X"4E",X"50",X"06",X"06",X"37",X"2A",X"06",X"37",X"2A",X"AA",X"A4",X"37",X"20",X"C2",X"79",X"85",
		X"AF",X"86",X"B0",X"84",X"B1",X"60",X"A2",X"15",X"24",X"5D",X"70",X"0A",X"A2",X"05",X"A5",X"5D",
		X"29",X"0F",X"D0",X"02",X"A2",X"50",X"F8",X"8A",X"18",X"65",X"A4",X"85",X"A4",X"A5",X"A5",X"69",
		X"00",X"85",X"A5",X"D8",X"60",X"A2",X"0C",X"A9",X"00",X"85",X"8F",X"8A",X"4A",X"A8",X"B9",X"8D",
		X"76",X"C5",X"56",X"90",X"70",X"86",X"3A",X"20",X"2F",X"76",X"E0",X"0C",X"D0",X"03",X"18",X"65",
		X"3D",X"20",X"BF",X"76",X"86",X"19",X"84",X"1A",X"A6",X"3A",X"E8",X"20",X"2F",X"76",X"CA",X"E0",
		X"0C",X"D0",X"03",X"18",X"65",X"3F",X"20",X"BF",X"76",X"86",X"1B",X"84",X"1C",X"98",X"10",X"0B",
		X"49",X"FF",X"A8",X"8A",X"49",X"FF",X"AA",X"E8",X"D0",X"01",X"C8",X"C0",X"04",X"B0",X"3A",X"20",
		X"43",X"78",X"A0",X"00",X"A6",X"3A",X"E0",X"0C",X"D0",X"13",X"A5",X"56",X"29",X"07",X"0A",X"AA",
		X"BD",X"9E",X"4E",X"91",X"27",X"C8",X"BD",X"9F",X"4E",X"91",X"27",X"D0",X"13",X"20",X"2D",X"76",
		X"98",X"A4",X"37",X"91",X"27",X"C8",X"E8",X"20",X"2D",X"76",X"98",X"CA",X"A4",X"37",X"91",X"27",
		X"20",X"38",X"78",X"A6",X"3A",X"CA",X"CA",X"10",X"82",X"A5",X"56",X"49",X"7F",X"C9",X"40",X"90",
		X"0B",X"4A",X"4A",X"4A",X"09",X"08",X"AA",X"A9",X"20",X"4C",X"53",X"79",X"60",X"84",X"37",X"A5",
		X"91",X"F0",X"1B",X"C9",X"02",X"90",X"10",X"F0",X"07",X"BD",X"7F",X"76",X"BC",X"10",X"4F",X"60",
		X"BD",X"71",X"76",X"BC",X"04",X"4F",X"60",X"BD",X"63",X"76",X"BC",X"F8",X"4E",X"60",X"BD",X"55",
		X"76",X"BC",X"EC",X"4E",X"60",X"00",X"FE",X"FF",X"FF",X"FE",X"00",X"FF",X"00",X"00",X"02",X"02",
		X"FF",X"00",X"03",X"02",X"01",X"00",X"01",X"FC",X"01",X"FF",X"FF",X"02",X"00",X"00",X"FF",X"00",
		X"02",X"FF",X"00",X"FD",X"00",X"01",X"00",X"FF",X"FF",X"00",X"FF",X"03",X"00",X"00",X"03",X"01",
		X"FF",X"FB",X"00",X"01",X"FF",X"03",X"01",X"FF",X"FD",X"01",X"01",X"00",X"03",X"5D",X"60",X"64",
		X"6D",X"70",X"74",X"7F",X"A5",X"61",X"4A",X"4A",X"4A",X"C9",X"08",X"90",X"02",X"A9",X"07",X"85",
		X"3F",X"A5",X"5F",X"4A",X"4A",X"C9",X"08",X"90",X"02",X"A9",X"07",X"24",X"5A",X"30",X"05",X"49",
		X"FF",X"18",X"69",X"01",X"85",X"3D",X"A5",X"74",X"4A",X"4A",X"29",X"03",X"85",X"91",X"60",X"A0",
		X"00",X"85",X"38",X"0A",X"A5",X"56",X"85",X"37",X"90",X"02",X"A0",X"FF",X"84",X"39",X"A2",X"00",
		X"A0",X"00",X"46",X"37",X"B0",X"03",X"D0",X"0A",X"60",X"18",X"8A",X"65",X"38",X"AA",X"98",X"65",
		X"39",X"A8",X"06",X"38",X"26",X"39",X"4C",X"D2",X"76",X"00",X"32",X"5F",X"9A",X"B5",X"CD",X"EE",
		X"FB",X"FF",X"00",X"80",X"C0",X"40",X"00",X"02",X"05",X"08",X"0B",X"0D",X"0F",X"10",X"11",X"12",
		X"13",X"14",X"16",X"18",X"1A",X"1C",X"FF",X"EE",X"0C",X"EB",X"08",X"EA",X"04",X"E9",X"FF",X"EA",
		X"FB",X"EB",X"F8",X"ED",X"F3",X"F1",X"F0",X"F5",X"EE",X"F8",X"EB",X"F8",X"00",X"F9",X"FD",X"F9",
		X"FC",X"FA",X"FB",X"F8",X"00",X"F8",X"FF",X"F8",X"FD",X"F9",X"FC",X"F8",X"00",X"F9",X"FE",X"F9",
		X"FD",X"FA",X"FC",X"F8",X"00",X"F8",X"FF",X"F4",X"12",X"F1",X"10",X"ED",X"0D",X"EB",X"08",X"EA",
		X"05",X"E9",X"01",X"EA",X"FC",X"EB",X"F8",X"EE",X"F5",X"F0",X"F1",X"F2",X"EE",X"F8",X"EA",X"FB",
		X"EA",X"FD",X"EA",X"ED",X"F3",X"F1",X"F0",X"F7",X"EE",X"F8",X"EB",X"FD",X"EA",X"03",X"EA",X"05",
		X"EA",X"08",X"EA",X"04",X"EE",X"FC",X"F9",X"FD",X"F8",X"FF",X"F8",X"01",X"F8",X"FC",X"FA",X"FD",
		X"F9",X"FE",X"F9",X"00",X"F7",X"01",X"F8",X"FD",X"F8",X"F9",X"FC",X"F9",X"FA",X"FB",X"FA",X"FC",
		X"F9",X"FD",X"F9",X"EA",X"FC",X"EB",X"F8",X"03",X"F9",X"04",X"F9",X"05",X"F9",X"06",X"FB",X"FB",
		X"EA",X"FD",X"EA",X"03",X"EA",X"08",X"EB",X"0C",X"EE",X"0F",X"F0",X"13",X"F3",X"15",X"F8",X"16",
		X"FB",X"17",X"FF",X"16",X"04",X"10",X"F1",X"12",X"F4",X"15",X"F8",X"16",X"FC",X"03",X"F9",X"04",
		X"F9",X"05",X"FA",X"07",X"FA",X"07",X"FC",X"02",X"F8",X"FF",X"F8",X"00",X"F7",X"02",X"F9",X"03",
		X"F9",X"04",X"FA",X"FF",X"F8",X"01",X"F8",X"08",X"FE",X"08",X"FF",X"08",X"00",X"07",X"02",X"07",
		X"FC",X"07",X"FD",X"08",X"00",X"08",X"01",X"0C",X"EE",X"0F",X"F0",X"13",X"F3",X"15",X"F8",X"16",
		X"FB",X"17",X"FF",X"16",X"04",X"15",X"08",X"12",X"F4",X"15",X"F8",X"16",X"FC",X"17",X"01",X"16",
		X"05",X"15",X"08",X"13",X"0D",X"0F",X"10",X"0B",X"12",X"08",X"FF",X"08",X"00",X"06",X"FC",X"07");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
