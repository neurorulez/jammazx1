-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D7A959F33CC4F679896798953D1E52716A664EC193324442C9000009B232165F";
    attribute INIT_01 of inst : label is "2EF1226F122EF1226F122EF3091248B244922C91248B245922C91248B24492A4";
    attribute INIT_02 of inst : label is "DFF1659B3743E51E13074143122EF1226F122EF1226F40D8CE338CE321226F12";
    attribute INIT_03 of inst : label is "F69FE27E33FF19ECA2766CA36423F4236425642564295AC6B162BB06185CCBF0";
    attribute INIT_04 of inst : label is "A450B2164C414B210B28CB66CB1642167774244FB53ECD29E431F421F50FA455";
    attribute INIT_05 of inst : label is "5E9264916489E06DB86B05EAD06047D080A5530082954C0A0A4D30182934C020";
    attribute INIT_06 of inst : label is "AF5A48F1A28410416D6F79C9CDB12F625EC04BDA897B10D526BF8D5F01AFEA32";
    attribute INIT_07 of inst : label is "15B33E4988D12C7669999A7493268D07511E767CD301A26C334EC684F70299B2";
    attribute INIT_08 of inst : label is "387996E23E5B88F9F18FA0E33EBC47D9B400ECEE7307A5CC96FD6FD266EFF7CD";
    attribute INIT_09 of inst : label is "69A1AB7C4A4DB051A85EE424BCE869F527518EB4257C49FB2268F34FFA4CC113";
    attribute INIT_0A of inst : label is "A3477CEF9DF3BE77CEBD2814A052814A052814A052814A052814A04EA4C1FFEF";
    attribute INIT_0B of inst : label is "CD4611B23CD0D4AE0330703B2223604C15525521074E465897606C7A3D1E8F47";
    attribute INIT_0C of inst : label is "0000000BCE51B187EF2C35979E73BFF8A80FC4BDE72815B0DCDB19A236E7AB5A";
    attribute INIT_0D of inst : label is "2F9FEBF85210E5BAB796EADE56F2B7956F2ADE5BCB6BBBB95654DAD000000000";
    attribute INIT_0E of inst : label is "4EBCEB6A0BD31CF9D79EB801550366489D9F9820035507D0FAFB3D73CE3BD1BD";
    attribute INIT_0F of inst : label is "24924924924927D55D37B3B5CCCDF3FBBB9D7F4F4C3AF3D969052D634AA0BE7E";
    attribute INIT_10 of inst : label is "5BF3C67FEFE6D6947E928FD9A18E77CD3E7A4FFFFFDDBB9B99DDDBBFDDFF30C9";
    attribute INIT_11 of inst : label is "56DE85BD0EF5921BD840F7FC67AAD79E4BF35FF3811441FE4129EDC48939B30D";
    attribute INIT_12 of inst : label is "C85243B25492E493B12B66F1B4FC4EC3FFF3722FD69EE65FED2D00B52B58D62C";
    attribute INIT_13 of inst : label is "164964964964964F5559E4BFDE6B84AB35492AC9524AB35F92EC2626BF5D237C";
    attribute INIT_14 of inst : label is "61989D060B07FD699B9D0683442766FB6F37B117EF79751326DED69C9B96B937";
    attribute INIT_15 of inst : label is "EFF8D3980D24E2DE73ED9C8F365CF301A6DBF390FB30FB2403937714143F989D";
    attribute INIT_16 of inst : label is "84D7493D7AFBD0996EBBA4A2A96EB0D889716226FBCF799DBD0B7A1DEBC37B21";
    attribute INIT_17 of inst : label is "522753382EFBA3C7892D93C78F125B278F1E24B64F1E3C496C96F2F870D683A0";
    attribute INIT_18 of inst : label is "9834F860DC1A7C30660D3E183746BF0C19A35F860DD1AFC306798D1C061D7727";
    attribute INIT_19 of inst : label is "77D5AC6F56FB5DEDAA03D7FB77E351DDFFECFFF768D7E30668D7E183746BF0C1";
    attribute INIT_1A of inst : label is "AB65463B6CA3AC70CEA392E8E2DB72B13FADBC93FED6F5FB54A5BACEF4DACFD9";
    attribute INIT_1B of inst : label is "9676F841460B54019B88D701CEA3536D944490A4B9DCB645CEB4289A3EA38D1C";
    attribute INIT_1C of inst : label is "11663B19620000E8080E0080E8000E0000E8000E0100E8100E0100E8100E63B1";
    attribute INIT_1D of inst : label is "B0D62D6328001B10CBAA8F1DDA20BA81511110AAAAAAA5555556AADC3BFA1812";
    attribute INIT_1E of inst : label is "7454A8A9D1544EEEEEEEEC4ED531473142D13AFD556458A32A08B144C47119A5";
    attribute INIT_1F of inst : label is "6A2AF455A8ABD156A2AF455A8ABD153A2A7454A8A9D152A2A7454A8A9D152A2A";
    attribute INIT_20 of inst : label is "31F9239C255055F353EBC65B9F984F6216375D25F79D769F3DA2AF455A8ABD15";
    attribute INIT_21 of inst : label is "F3713CE984FBF0D3C40931C4FE27FF1AF57F3ABF9C464458574FE20235103A61";
    attribute INIT_22 of inst : label is "6311B11B69081245557E04021F52B58D62C54AF00E7AF40E7AF40E7CD44F9A09";
    attribute INIT_23 of inst : label is "79E300022C18001161FFFFFA204AAAB6A4EAF0EAF14A9098909890989B9B9B9B";
    attribute INIT_24 of inst : label is "6A8940599A0A84AAC994E4C8F131002C008588CA3F264C500B002162320FD805";
    attribute INIT_25 of inst : label is "592C964CCC04A55840E89695550A04260BE11179645D91658C17D56BD84FCB53";
    attribute INIT_26 of inst : label is "20D5D16465597D96D97EA0BA6B685B10048B798B5789282ACD3B2592C90864B2";
    attribute INIT_27 of inst : label is "8A01CD8AFAC4FA71DC567E59FD94CC3475ABDCE074E2EB0FACF8719BBC2E76A3";
    attribute INIT_28 of inst : label is "1C4466388834E1E9DC243B9212A24560D980202052C1961504D20706D86C0104";
    attribute INIT_29 of inst : label is "2D591125E5E5E584872F2F2F2ED6D4E8C58B31662CC598B3BEFBEFB6294FCC33";
    attribute INIT_2A of inst : label is "A157B9EE7E7B9A02D20C63181797889F06A455AABBC8AF0A458109F0302ABBB2";
    attribute INIT_2B of inst : label is "418C295185AA30A54616A8C295185AA30A54616A8C46231188C46231131189AD";
    attribute INIT_2C of inst : label is "5602F50ABE7CF9F3E7CF9F3F3E7CF9F3E7CF9DCF77BBDFC2FD579123F94B8651";
    attribute INIT_2D of inst : label is "1F5C02D7F63609C9C690326997F79EBDDEF610CFB0867B2BF968812A93ADED6F";
    attribute INIT_2E of inst : label is "B3A2B31C7456479164FFC8A86EB495220A2C6090A77A1A7C98368D1515281B1A";
    attribute INIT_2F of inst : label is "22AB1A7409BA49A0801A40F1D9591C765647B3B2B31C745647B3B2B31E745647";
    attribute INIT_30 of inst : label is "6DD3DD5BB4C2B0C5A006D2A2E84F2A6EE581671DA356E6E6E2F2F6BECFECCD8A";
    attribute INIT_31 of inst : label is "A4CDAFF0CE41208148A212BA87476DB642924924924924924D31094EF2690AD1";
    attribute INIT_32 of inst : label is "3790B79358043D1633189E976353D8EADFE6B7FED1A0031C600C20A95AC6B162";
    attribute INIT_33 of inst : label is "2144000C71C070BE1C3705A8000638E028412210018E380A104AC000C7180708";
    attribute INIT_34 of inst : label is "4B8522D5676356167AA88F50000C718030B60C170490B2009379F9882B5BC16F";
    attribute INIT_35 of inst : label is "6AA379A002A0F4D191AD5DE5811A8EF6774B89CCB065A9607682A4479B53B3E7";
    attribute INIT_36 of inst : label is "CA6B948963C66985A65913A9CADC3A78D202CDC2BA0E542C4C84C1A6A531387F";
    attribute INIT_37 of inst : label is "66D5EAC57852393FDFEFFDDDDB091AE96A029169A7A14905E8248AF013457808";
    attribute INIT_38 of inst : label is "800A0016152B175D252C962EBA6B474EA7CC520E55343D73A4CDD12AE4D51515";
    attribute INIT_39 of inst : label is "AC9209276490492B248249D92412460400E1860049009001282BC310F8078005";
    attribute INIT_3A of inst : label is "13398362203A3A9061ABBFC738B02602D802C9309236498490B24C248D926124";
    attribute INIT_3B of inst : label is "05D7422360E029E55ABBCE0525E648A5291809C3504F781F2A0B00761014C406";
    attribute INIT_3C of inst : label is "53CD115456624F9E8DE156F7AC685D0336D22DB698041823AAAAB8A88CECD895";
    attribute INIT_3D of inst : label is "80210040000288000004210801C0210840000000A0008021080045515B57B0A9";
    attribute INIT_3E of inst : label is "1004010000020008001084200310000000020000800000802100420070080210";
    attribute INIT_3F of inst : label is "58D24D49A93526A4D49A93526A4D49A9E53CE993CEDB279C9E56CF38C0200002";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "6C43800BBED8477DB077DB0591A48CF61F261FC98635CB10950000418E48848C";
    attribute INIT_01 of inst : label is "00DE500DE508DE508DE500D9B285940CA0650B285940CA1650B285940CA0658B";
    attribute INIT_02 of inst : label is "0E828A24C889B74F311232E5E508DE508DE500DE500DD97D0741D0740E508DE5";
    attribute INIT_03 of inst : label is "063FE9AC8D6F4E93E5E3490A008A908A008E008E00F2500532A52B2ED8FF89F4";
    attribute INIT_04 of inst : label is "7E056C4034B31284424210109084888482882898C00A7B62D898D898D846D0BB";
    attribute INIT_05 of inst : label is "B845022A11400FC0C7C033078E9EBC543F7F3EB65968B3F5F7EBEB45968B3F5F";
    attribute INIT_06 of inst : label is "F8F1278B047F6FF6D658851E580EDC0DB059B709B6C1272C1B6036E166DC25CC";
    attribute INIT_07 of inst : label is "356CE0F25122ECF9962A6DC36ED970169AF089C1A4F645FCCDB819AB1849CD25";
    attribute INIT_08 of inst : label is "26C42D316CB445940F7805306DB20CBB4A7949114CEC7B1FB23622459202FFD8";
    attribute INIT_09 of inst : label is "C41E5803D9D844675BF0985DE1109B114022344BDB81B60B35B40DB902A8BBBA";
    attribute INIT_0A of inst : label is "FC640981102604409815997665D997665D997665D997665D997665BDFBB30078";
    attribute INIT_0B of inst : label is "9DFFFB4672792009F7BA8F73B48F64ECBDA4F7626DDB5B39BFE4C58FC763F1D8";
    attribute INIT_0C of inst : label is "FFEAAA823882CA391C44CA3AF434400178277970186AA33386672459800C2FFB";
    attribute INIT_0D of inst : label is "560FEFFB3B3B10B4A842D2A1050828415082A1042091504554F17C000005555F";
    attribute INIT_0E of inst : label is "192105E6A59A696B242059921E658C31E4C420913C1E6BDF6F5C45B1025CA61A";
    attribute INIT_0F of inst : label is "184184184184191577C955C6C48525AFAA67971669E48429B769B6A5BBCD54B4";
    attribute INIT_10 of inst : label is "E123C9F81C0D48B1121E236B55DFFD5A60D487FFFE00000002464442222F0404";
    attribute INIT_11 of inst : label is "A039147321CC67073F9ACFFDB351D1619609A80C223923FE92C70133664448DA";
    attribute INIT_12 of inst : label is "23811508E847036C46DCAD04093C8CB89D0885882D3109105A055C0E4A00A654";
    attribute INIT_13 of inst : label is "8820C30820C30822A304196030BE7B40CF065936E1B62DB065888BC1D6804951";
    attribute INIT_14 of inst : label is "B3E6339B3D8FF3B3E5339B3599C81D0C02CA424400A29E448F295B3BB45EF768";
    attribute INIT_15 of inst : label is "9FFB6310581BE785ED977B261C9B200B036704627002701607768F61297FE633";
    attribute INIT_16 of inst : label is "494DC25DCF5C752A976FC956F4900149140224558DD8BA107228E64398E0E7F5";
    attribute INIT_17 of inst : label is "C9ECC8F5A084F54AD412A56A95A8254AD52B504A95AA56A0952BABA899490459";
    attribute INIT_18 of inst : label is "43C9115AA1E488AD58F24456AC39022B541C8115AA0E408AD587CF224F238CEC";
    attribute INIT_19 of inst : label is "868A28BE68D457D155F608AFA07CBD12DFF92FF58F244AD58F24456AC79222B5";
    attribute INIT_1A of inst : label is "C2266607C4C05A6B030042F014F47FC280036A0600F8E073F14A201F891B20CB";
    attribute INIT_1B of inst : label is "C31E7000801D2801534006906D80353C24A04948D34CA242AF1200D550D04C02";
    attribute INIT_1C of inst : label is "4218319C348080E0080E0000E8080E8000E0000E0180E8100E8180E0100EC319";
    attribute INIT_1D of inst : label is "6BCD1A96F7F7ADAD7F3E5C3E73BDE340EBEBEA19999999999998CC4C94B55C7F";
    attribute INIT_1E of inst : label is "E89BD13722614BEBEBEBEBE12BEC8842BF624F5AA238A59086714B303CBFF793";
    attribute INIT_1F of inst : label is "244C6898D131226244C6898D131226F44DE89BD137226E44DE89BD137226E44D";
    attribute INIT_20 of inst : label is "7B02CF5399A68E03F61E6BE2605C94C2D267EEFA165FB9F0B344C6898D131226";
    attribute INIT_21 of inst : label is "140A43B669060D2F3FBCA628014000A6CB80E5C073DA8BA489B014CF5E7FED9A";
    attribute INIT_22 of inst : label is "97A2FA2FF477B4289B81A914F0E4A00A654A3B0EFC830EFC830EFC850E90A152";
    attribute INIT_23 of inst : label is "B2F67528F9B3A157CB00000158BA49B7DB9CCF9CC8B96771277127713F3F3F24";
    attribute INIT_24 of inst : label is "A1582B3E00D4CD1D572FDFBBCFEF7D49954E1383A0FDFBCF52655384E068397F";
    attribute INIT_25 of inst : label is "3E1F0F81B3DFCFB3BEAD205A2EF7797F5CFCEFE2CFFB3FCE56EE625C4FA0FAEE";
    attribute INIT_26 of inst : label is "5FA622CFAAAC5A80AC51C5CD000E00FFFF65F3FC2CCBC79552F7C3E1F0F7F87C";
    attribute INIT_27 of inst : label is "1CFCF39759CA002F4EEF043C14FB85C8AB972FC5EFC936759E062F65C7F7EFCD";
    attribute INIT_28 of inst : label is "239AFC4F745D5F52534BCA256FFFEECB9F15B5B503971C9DA799503DF2F914AF";
    attribute INIT_29 of inst : label is "DFB3E2C323232329391919191B6B7A17CB97E2FC5F8BF134A28A28A697E8B77E";
    attribute INIT_2A of inst : label is "77E37FFEF7FFBD69E97084777E7E69002970EF31259116DD096A100149717767";
    attribute INIT_2B of inst : label is "2A5EA36BD46D7A9DAF53B5EA36BD46D7A9DAF53B5EAF57ABD5EAF57B3FEBDFDB";
    attribute INIT_2C of inst : label is "88700C75681020408102040408102040810201A0804021B7379E5FD8EBA18B33";
    attribute INIT_2D of inst : label is "F923703C1B49DA1A21293590E88659020108AC90456483C4400562EF6E73939C";
    attribute INIT_2E of inst : label is "AC44557B8A8A8EB73B002B13900EE1B4D4D5A74FA9976102FAB951A22633E435";
    attribute INIT_2F of inst : label is "4C44E54B5AB5BEA66E796F462A2A3B8A8A8EAC44557B888A8EAC54557B8A8A8E";
    attribute INIT_30 of inst : label is "B6762339EC94414E9B5E40440D6FD49D523806DA64C9C9C9CDCDCD49CC9CC3E5";
    attribute INIT_31 of inst : label is "2FF4F43DF188C413275B79F3FE7BB6DB6D6186186186186183BC77CD14F3271A";
    attribute INIT_32 of inst : label is "CD2D4D2E93333F3ED5299FDAA533F3454FE554FEAB0554E30BF7E772500532A5";
    attribute INIT_33 of inst : label is "5A9C15538C2AFFBEBFEF3AFDAAA9C6157ACEB77AAA718DFBF3AF955538C6AF59";
    attribute INIT_34 of inst : label is "B22BB7DF39B4CBABFD913FD6D5538C6ABFB6AFCF39A586E5A6D3F8265A26A29A";
    attribute INIT_35 of inst : label is "84C692DA251E0AABED7892C96A2B6D69B4D5D1B9DB8AD2BF6C3536B9661C4418";
    attribute INIT_36 of inst : label is "9DA4AD72ED9C36BA7565EE76B92EED952175456520DDA678BBABBF70D2A6A745";
    attribute INIT_37 of inst : label is "2DE60788B6E877807038066237E8A912673B4A57BD3FB0B2994F5948A6ACA452";
    attribute INIT_38 of inst : label is "722CE45B52D15AD6CE05A2B5AD9C0EDDA2556DF4D64ED0CDD90232EB0B266222";
    attribute INIT_39 of inst : label is "3B089C13D84CE09EC227047613382FDAD5DADFF22EE45DC8B2A5B4B2656B7916";
    attribute INIT_3A of inst : label is "54E75E445DD94D6AABD44FCCC14748E873FBB089C17D84CE0BEC227057613382";
    attribute INIT_3B of inst : label is "2A206D457DBD1AEDE12595FE0DFCADEF7A0665E08CD7FAE214722EF45E8D0BBA";
    attribute INIT_3C of inst : label is "2816A2668525A0657B52F5ED6B916E254DB85B6D925CC1C4547441F1D3130B6A";
    attribute INIT_3D of inst : label is "0401004000840802008020004284010040100021020080200042499A11A345F7";
    attribute INIT_3E of inst : label is "10040100021C2008020080010C00802008020087080200802008001081004010";
    attribute INIT_3F of inst : label is "A5B8000000000000000000000000000000001A40013C8002000400C784010040";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "AA4A80EA288624510C451084702BBA955D521A848690CC5000000004A6628484";
    attribute INIT_01 of inst : label is "82A7D82A7D8AA7D8AA7D8AA23EE1F60FB87D8BEE5F62EB87DCBEC5F72FB17503";
    attribute INIT_02 of inst : label is "1A3028F162D9A705100550A67D8AA7D8AA7D8AA7D8AA1180401004010FD82A7D";
    attribute INIT_03 of inst : label is "94954B54B6AADB766307522A002A902A002A902E00508E142C28420AD26FA09E";
    attribute INIT_04 of inst : label is "4994481080E55241548A365122A902A009DC9DF7195924A8002A902A9150042E";
    attribute INIT_05 of inst : label is "A17D9BEC9F66EEA5DEA10E834CECEA043249B6936DB6924DB6D24DA4924DB692";
    attribute INIT_06 of inst : label is "54A8C94283CDA6937D747A64D4BFD4AFA149F4293EA533AA5F50BEA127D4271F";
    attribute INIT_07 of inst : label is "10D35259B3D3A863D400F50BAA1D50B4D3A8E6A4B323A7681EA04ECEEF40DD49";
    attribute INIT_08 of inst : label is "B0A49A411269044B6A54E0C0132822629E60EDCC330A50EA569269276634CB14";
    attribute INIT_09 of inst : label is "A1AF543A82837B7A90A8666151CCC2856733B77DEA15D52A17F70EA172E6C2A9";
    attribute INIT_0A of inst : label is "A5CB746E8DD5BAB746EF6E9DBA76E9DBA76E9DBA76E9DBA76E9DBA60BE61FFD4";
    attribute INIT_0B of inst : label is "50A522726CD3D28632A8E32A33744088693BA5D38A74DC90A840A6BA5D2ED76B";
    attribute INIT_0C of inst : label is "84411DD7CF7337CFE7BCF7CD2BA73828501B7F50EF4381A14992732636CA0425";
    attribute INIT_0D of inst : label is "571D53549C9C65A60D96983651B28D941B283656CAEFAED803764AE77BAEE208";
    attribute INIT_0E of inst : label is "2C964FD330E79E9592CAF419638F603871D140C18F639D5F65B67A784596D41D";
    attribute INIT_0F of inst : label is "20828A20828A23001F6DFF61C2007A4ABF72ED1B9E325970EE9E1DCF7473EF48";
    attribute INIT_10 of inst : label is "B2DE9B07E1AA1A55490AA92281D73A1451A083249357555755311131315A188A";
    attribute INIT_11 of inst : label is "0E94152824A154529F50A6A9D39A8509D52EE277A25C5354C38C20CCDC733714";
    attribute INIT_12 of inst : label is "BEE9F64FB37D93AA17502A7591C082B162603B226A28764494885C4A11C28585";
    attribute INIT_13 of inst : label is "145104104145145635429D509A6B3D72EA97543EA1F42FA17D40AB536D110B05";
    attribute INIT_14 of inst : label is "EEB2B8CEE70AA8EEB2B8CEE715A95A719CAD93112CD9A333AC364E9629B5AC53";
    attribute INIT_15 of inst : label is "4D53AA581424C54651C994C627540102849377A0D480D00142C532D71DD532B8";
    attribute INIT_16 of inst : label is "9FC5C7F745B6DBFDFE2F9FE2F9FAA11CC542731243D47B51292A5049420253C1";
    attribute INIT_17 of inst : label is "134B1359BB39A7AF5C3FFFAF5E387FFF1EBD70FFFEBD78E1FFFD6D68C9DFC649";
    attribute INIT_18 of inst : label is "E8ED593E6476AC9F3A3B564F995D8B27CCAEC593E75762C9F32D070C470DB34B";
    attribute INIT_19 of inst : label is "C9DE5DD3393CBA72080280295556C4BF754FBAA6CBB169F32BB164F9D5D8B27C";
    attribute INIT_1A of inst : label is "E9D74E493AE4952AD0D48629213C8D436C6D8C8479290D84A96C46D04DA39B73";
    attribute INIT_1B of inst : label is "EB9D1800420E70016141028205042AB2FC3F8D27E9219DCEC282A6D096E49D24";
    attribute INIT_1C of inst : label is "1472658EB18180F8100F8180F0100F0180F0100F8100F0100F0180F0180F6658";
    attribute INIT_1D of inst : label is "078081CC67463B31D2B0D4582A656B8014015507878781E1E1E0F0109EBF444E";
    attribute INIT_1E of inst : label is "8CDF19BE33754ABFEABFEAB7BF58CD6BD3B3E5B3F31F7CC9C33EF99A76472300";
    attribute INIT_1F of inst : label is "066E2CDC59B8B37166E0CDC19B8337C66F8CDF19BE337C66FACDF59BEB37D66F";
    attribute INIT_20 of inst : label is "AE9193B3BB7DF39AD336CE33AC90EBC270E659A335196699A866E0CDC19B8337";
    attribute INIT_21 of inst : label is "2313A43B0E95218282369F5C4AE26530A0B238591C3FCC38CDDC871AC6930EC3";
    attribute INIT_22 of inst : label is "4433833807BA3F3CDCE42E1729A11C28585084C08B4CC08B4CC08B48C0E9181D";
    attribute INIT_23 of inst : label is "FB1394287E9CA943F4B366C870EB2C2524CCA4CCA0E9D991D991D991C2C2C2D2";
    attribute INIT_24 of inst : label is "E6F0DE970B1F0FEF9831A346A0D1C16D15CF9D44991A34605B4573E7512644DE";
    attribute INIT_25 of inst : label is "0381C0E6ECCC7EFFE2CDBFDF30E4766457A0189BFA27E8EB18F9B378D19BC3DB";
    attribute INIT_26 of inst : label is "71FFB3EBF3E44A40A440656F7F25008CCFC71B163E5FE73F164870381C930E07";
    attribute INIT_27 of inst : label is "86F38439C81DB826BCB0DC0374CF7E6DEC18B9A19129BFFC81B236B71C5C9067";
    attribute INIT_28 of inst : label is "B4861B690C13C6FAA0D2D44141870BFA548D050771F48F95225277523E1F0C3F";
    attribute INIT_29 of inst : label is "E0FAF372525252181A92929290080A2E0C18DB1A636C69A5451451408EB0000D";
    attribute INIT_2A of inst : label is "93B8A12941421264A47AD76C450503892C58FA3BFEF99B56CDEB38996159CCFD";
    attribute INIT_2B of inst : label is "9F4A0B894171282E2505C4A0F8941F1283E2507C4A25128944A2512860694494";
    attribute INIT_2C of inst : label is "4D3037B9A72E5CB972E5CB9193264C993264C99E4F2790F59EF533C6B2DC0A17";
    attribute INIT_2D of inst : label is "A4323029F664D3130BF194DCCA7514793C9678E9B3C74BA65801C3AC933D49EA";
    attribute INIT_2E of inst : label is "C677EFA4CEFDE9837E99E39AD9B6D61F3EF3EF8E2CDC7ADEEADFE9C77331B67F";
    attribute INIT_2F of inst : label is "6EE72C205B3092CCE46367133BF7A4CCFDE9C677EFA4CCFDE9C667EFA4CCFDE9";
    attribute INIT_30 of inst : label is "D894896D3DDFE39F3E7061FF394A4EAE3318065D3264B4B4B4A4A4648A4AA98F";
    attribute INIT_31 of inst : label is "50A85A2585F4FA6DD9EE6DABB5726DB6CE38E38E38E38E38E633BAAC92683533";
    attribute INIT_32 of inst : label is "F1B171B2DA2229308A391481472290060D55A6AAB507D79EBBE3E7D08E142C28";
    attribute INIT_33 of inst : label is "62E6955E7AFE8DA1A3543C2A4FAF3D5F46CF4A93EBCF57D1B3D2C9F5E7AAFAF9";
    attribute INIT_34 of inst : label is "EB2E39181B370D2D5219EA1D155E7AEFCFA9F3F43E161726171B50B06138E2E3";
    attribute INIT_35 of inst : label is "CEE63FB2679DE67324D1FF7DEB33ACDCE2DFFD9F73F799E772C7C7CD574F718C";
    attribute INIT_36 of inst : label is "D6FF8C5A8B9A3F9B933DFC925FDEDFDEB11701B2DB17F86FF63F66D2E397992F";
    attribute INIT_37 of inst : label is "0CFF450CDAB63AD3C9E4E8889B303FFF490AD24EB9A7FCD3697669B0BB34D85D";
    attribute INIT_38 of inst : label is "1831306062187E4B6F01B0BC96DF164E9DDDB7BFE7724B67FD873B73ADB37773";
    attribute INIT_39 of inst : label is "51C6D4928E36A48471F524A38FA924148682141831306060C4C4243301084C18";
    attribute INIT_3A of inst : label is "56D6AD64E1F96853D69EEA35FE5973287D111C6D4908E36A49471F524238FA92";
    attribute INIT_3B of inst : label is "9FF7917AA9491B08A7FEFCCF081E8D08434E44098CFC50F3967B2486548D9C3E";
    attribute INIT_3C of inst : label is "76FBD7375C59DB7FCE78A779CEDE7BC7E92A52495274CEE7EF9FBEDEFBFBFB77";
    attribute INIT_3D of inst : label is "80200802100200401004010801802008020084008010040108019CDD74F8F91C";
    attribute INIT_3E of inst : label is "0080200840080100401004200410040100401003004010040100420040080200";
    attribute INIT_3F of inst : label is "319A244488911222444889112224448889114915149A2A28A895177B00200802";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "CE08802F75662EEAC8EEAC8E3032B2815C10284C0B81AD440600006D2D6A2014";
    attribute INIT_01 of inst : label is "CB791CBF91C3791C3F91C37F48C446223911C08C046033811C88E446223119C8";
    attribute INIT_02 of inst : label is "120138A142B74E58118050E791CBF91CB791CBF91CB715F8C2318C23091CBF91";
    attribute INIT_03 of inst : label is "839FE71874CFB2640766522200229022002290220058218AA8C1FDE47DD5CB94";
    attribute INIT_04 of inst : label is "4D904814B4D54281900C8064022002203A4D24D3115A042A1832003201101437";
    attribute INIT_05 of inst : label is "303989CC4E602AE15AE30582C4D6DE401269249B6D369349269B69B49A4934DB";
    attribute INIT_06 of inst : label is "FCD877CB80ED369B693CFA6EDC3918B2314A472948C534CE4672CCE5299CA6F3";
    attribute INIT_07 of inst : label is "09F3B30F05AB64AE662F99888E44729C7B7867661E0B568CF3310D2D3940D948";
    attribute INIT_08 of inst : label is "16E4B661BED986F9F39C21E1BECC37D5947824CD73663AE81400400764A4850C";
    attribute INIT_09 of inst : label is "6329980CF6F7FAFF9FF8E569F0CED39C7911936D3396672D566603311CEC59B3";
    attribute INIT_0A of inst : label is "65EBED7FAFB1FE3EC7FBF7EB56BF7EB56BF7EB56BF7EB56BF7EB56ED3E71501C";
    attribute INIT_0B of inst : label is "9E63713838A9B18E337A631DD66BE55CEC33B1D36E74ADF99FE666B75FAD97CB";
    attribute INIT_0C of inst : label is "85050A09E7DBF3CCF3EEF3CFA317F828621F447029610113CDFB7BF7DB76339D";
    attribute INIT_0D of inst : label is "14BFF5FD8585E537E794DF9E5CF2E797CF2F9E53CA7AFEBFFF47ADCA01414282";
    attribute INIT_0E of inst : label is "249E4336B669A49493CA2D5B6387761E3D80C4D9A7638DFFF92E6F69C7779215";
    attribute INIT_0F of inst : label is "69A61861869A6B7FCC2F332D87C3925EAAB48B99A692793CEE8E1D877471E24E";
    attribute INIT_10 of inst : label is "729D4BC375067114006280018A51860CB33C444926999BB99B99B99B9B955CDA";
    attribute INIT_11 of inst : label is "3B8DDB1ABC6D16B1AA576BFC9E96C72C47072914AB575BFE7B7EB5CDDF33778C";
    attribute INIT_12 of inst : label is "1C80E407213B00CE199C36179802FE995E6932A2461865448C7C246B04315518";
    attribute INIT_13 of inst : label is "B4D34D34D30C30C62D50C470CB49667223919888E447023011C26AE04BA10201";
    attribute INIT_14 of inst : label is "C879AFBC9EAC1FC878AFBC96E52A56311C298BD1189F93BC68267D4D594AFAB2";
    attribute INIT_15 of inst : label is "D7F932921CFEBFCA376D8DDD7BEDB0439FDA94B09010901DE1AB2A640F00F9AF";
    attribute INIT_16 of inst : label is "EDDDB968392AE9B0DAECE58CC65E69DF6CD37DA7EB4A68931BBE3778D2D6356A";
    attribute INIT_17 of inst : label is "6E9B6E85FB1FB2A54FCB16850A1F962D4A953F2C5A14287E58B5E0E468ADB36C";
    attribute INIT_18 of inst : label is "CA7C6A68F53E35347A9F1A9A390F8D4D1E87C6A68F43E3534738BC380A39F25B";
    attribute INIT_19 of inst : label is "D04686511A0D0A3457D5DD758E32F5CB3FE59FF2E9F5B347A9F5A9A3D4FAD4D1";
    attribute INIT_1A of inst : label is "C086425110C5303814250221420D225125B4C6A02A4A568927BE8B4A97C0C99A";
    attribute INIT_1B of inst : label is "D74C8000000C0401C1C1438287056072A4680880C39488438226568C24850428";
    attribute INIT_1C of inst : label is "0852638D70008060080600806008060080600806008060080600006000066638";
    attribute INIT_1D of inst : label is "9312A5F5C7E7FEBFB3565E4E337EE1C0155400007F807E01FE0300DEEF6E9DE2";
    attribute INIT_1E of inst : label is "17662ECC5D154AAABFFFEAACE7BC4631BCB5792F91567F59CD6CFEB26AEEEE24";
    attribute INIT_1F of inst : label is "5BA295452ECA5594AB297452E8A5D99AB337466ACCD599BB315662E8C5518AA3";
    attribute INIT_20 of inst : label is "4790D1501B7DF795F3AE959D4C9ED0D79063D963AF4F65997BAA2B7656A8AD51";
    attribute INIT_21 of inst : label is "2D93F42F4FD5A8AFA32C71244923651FEA32951D4E066435657CA68BDE5B0BD3";
    attribute INIT_22 of inst : label is "6463C634373F722C766525538DB04315518383608ECB608ECB448FEB40D9681B";
    attribute INIT_23 of inst : label is "EB1B23A4E5DD1D273E72E5E96CF9458766C9EEE9FDFBB399B399BBD9E3A3A3FA";
    attribute INIT_24 of inst : label is "E35048BB8B0709A1A85362C278B2056451FB1E437D162C8159147EC790DE427C";
    attribute INIT_25 of inst : label is "2592C96222832CC8F25CB68F18F9495946A53835300C8030D7BBD1B48BED85A9";
    attribute INIT_26 of inst : label is "39511120D2C6C06806C3346A4927A02B69E2AAFF122C67D6045CB2592C45964B";
    attribute INIT_27 of inst : label is "E579162EA916DA1DD6F96A25AC3EE9BDCE4C117F3968A99892DC1DDE4AF9B923";
    attribute INIT_28 of inst : label is "9FF19637A36CE58B25756495DDCE8B34F1F7DFD69C49E37BF8F769E70986EEF1";
    attribute INIT_29 of inst : label is "724C31B1939193AEAC8C9C9C8CEEAF7F060CB19732E65CEE49249249DE326BCB";
    attribute INIT_2A of inst : label is "573919E77A719F7D7CDC725E6363E0ED25B1B60ED758898746878E913918D990";
    attribute INIT_2B of inst : label is "8BE7BABDF7579EEAF7DD5E7BABDF7579EEAF7DD5EFF3FBFCFE7F7FBFBABCFD59";
    attribute INIT_2C of inst : label is "8F70233FB3264C993264C99D9B366CD9B366CCFF4FA7DA61CCFF7B7B10EC65F2";
    attribute INIT_2D of inst : label is "DE38F0196674410199EFAB788A5F7FFD3EDF3779F9FAE9477005B3E59B2BDD5F";
    attribute INIT_2E of inst : label is "8AAA331D554447ABCF9D70897ED7F613273A5D8FDD4F936DE5D0EAF11577DE27";
    attribute INIT_2F of inst : label is "A22289CB47176D5CFD6FFF1555191D5544478AAA231D5746478AAA331D574447";
    attribute INIT_30 of inst : label is "DDEEDEB98A6737DDBEBC4133B90F76A523B803AA1428E8E8F9F9EC44FC4DEAAA";
    attribute INIT_31 of inst : label is "EA09921AB764B249936E79B5F6BF4D34CE59659659659659631B3FD59BCB3BB2";
    attribute INIT_32 of inst : label is "60C560C4CE777A25AA93BD3552F7A6B297F9A2FF303736292C8B9DD8218AA8C1";
    attribute INIT_33 of inst : label is "8AC25458A4A20471C39EED306E6C5251073B0C1B9B149445CEC30DCD8A4B22E7";
    attribute INIT_34 of inst : label is "4D1F50CBB8EE042C74088EC4D458A4B20471C39EED191C3D1C0CA8CDC19054C1";
    attribute INIT_35 of inst : label is "EA3EE89BB79FF5C94FB36BAE8715D70D0A2718E606C6179E2EC9C2579936A2D5";
    attribute INIT_36 of inst : label is "92ED095F1B562F2B5E8B3148EB58BBCBB03604949B023846EC0EDDB871F176FA";
    attribute INIT_37 of inst : label is "9C9143044C3B1592A956BDFDE1509B4BD39EEAED185F7AA2D929516895A8BC4E";
    attribute INIT_38 of inst : label is "9B7736EDEF1CE669611339CCD2C2338516EA979A81A91926BDC31980B6F51111";
    attribute INIT_39 of inst : label is "8ECACEDC765676F3B2B3B79D959DB9BCC737999BB7376C6EDECE4767919C8DBB";
    attribute INIT_3A of inst : label is "67BDDB2635657E7AE7D7602DAC322F46CF9DECADEDEF656F6F7B2B7B73D95BDB";
    attribute INIT_3B of inst : label is "DB55D573BFDFD39E72D75CC9100366C6B0CCF719ED8E7FB9E7592FC25FA9C6AC";
    attribute INIT_3C of inst : label is "5B6FD19B8CB76DDBF6BCAB18C77CB39E7EF17DF6CB76EDA2B3B7AC1C1ECE93D9";
    attribute INIT_3D of inst : label is "39CE739CA6133184A508C6300188425294A108849CE5294A7201846E369D37EF";
    attribute INIT_3E of inst : label is "6738C63088CDC612942339C8442129C633942233339C6318CE508C044A5294E7";
    attribute INIT_3F of inst : label is "79DA224448891122244488911222444A995B4F1125D7234E8911B14F094A1084";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "0C3288CA08083000104101018EA8EC9E105B022EC0D1899040000006AC4C8693";
    attribute INIT_01 of inst : label is "CC9C1CC1C1CC1C1CC9C1CC99A4C7273939C98E4E7263939C9864E3261938C9C6";
    attribute INIT_02 of inst : label is "2ACA49224591A774A9D59AC5C1C49C1C49C1C41C1C41D172A4A02A0A0C1CC9C1";
    attribute INIT_03 of inst : label is "453555415E0A2F23140B044AB2C86AC8B2CA22CA2282C7D1C2A508374099AE84";
    attribute INIT_04 of inst : label is "0425116070B281D6D1121A9044A22CA210CF0CD46A4532523ADA22DA225102BA";
    attribute INIT_05 of inst : label is "30E94F4A7A5188167014B05420B0B16601248209041040048009040049209241";
    attribute INIT_06 of inst : label is "420510205636496DA682493402CC18D8318B0731E0E6264E706360E62C18C588";
    attribute INIT_07 of inst : label is "A1058996D572CAA12634418E0E72635182C40B132DBAE5828831EB4BDC6DEC10";
    attribute INIT_08 of inst : label is "2410E100658401940842970064002C88525D5019464108332A1AA0849A082912";
    attribute INIT_09 of inst : label is "96CC1CE212800E2C50848E4C0818984D6C333771830B071017073830C2C49001";
    attribute INIT_0A of inst : label is "92549A93522A4549A9348912245AB56AD48912245AB56AD489122400380A5512";
    attribute INIT_0B of inst : label is "008840CC266F6948A4820A4025D8178A8AAE2A02C9838B15A116124924904824";
    attribute INIT_0C of inst : label is "000040032C824B2D9640CB2C6806252D7EBB5073CC724AAB276C6EDDCD810484";
    attribute INIT_0D of inst : label is "476D4F5323231A2744489D11A889446A889511A224511046A881361084000800";
    attribute INIT_0E of inst : label is "2DB4420424DB6DBDB68A21929B76BA1BB6C60499369B6E8805826A30C482E75E";
    attribute INIT_0F of inst : label is "4D34D34D3451442A982D776AC94736E5403AE09B6DB6D134D26DDA46936D86DA";
    attribute INIT_10 of inst : label is "164C2D0496216129046D21A85B14A40208C2032491002002020220002240CC13";
    attribute INIT_11 of inst : label is "A1739AE73399E58E639C9AAAD8597119271C78E63A23235532D2411932064CC2";
    attribute INIT_12 of inst : label is "F4C7AE3D30E9860E2C1841466000D1150180CDC181059B8302EE45A058FA3854";
    attribute INIT_13 of inst : label is "A69A69A69A69A698B283927341B4F261838C1C64E3261830C9878C8021360D15";
    attribute INIT_14 of inst : label is "BEEA35DBEDAAA5BEEA35DBE5F9CD9146B2DC82E0A2C7A2ED8FB35BC304F58609";
    attribute INIT_15 of inst : label is "3555AE27425B35258DB66377D98310E84B6C472B510B511D94609EBAB1D56A35";
    attribute INIT_16 of inst : label is "ADBBFB7F458675BADDDF6DDDF6D99983B3330ED385D1BB26E735CE673BB1CC79";
    attribute INIT_17 of inst : label is "25912599CA88D72E5A5B372E5CB4B66E1C38696CDC3870D2D9B8282EC9ADE64D";
    attribute INIT_18 of inst : label is "8D7B653846BDB29C235ED94E15AF6CA70AD7B653856BDB29C22610A7A8A791D1";
    attribute INIT_19 of inst : label is "D8C6CC531B1D9A7677FFFF669292709B754DBAA6D5ED89C2B5ED94E15AF6CA70";
    attribute INIT_1A of inst : label is "0E102C96C2094B0125195592571D95436C6DEF272B2B2D8CA927C6D564E19B36";
    attribute INIT_1B of inst : label is "08033F7FFFE32C02380A5014E0A91E8C0993404730E121A969108015605959CA";
    attribute INIT_1C of inst : label is "4E08040080810008100081000810008100081000810008100081000810008040";
    attribute INIT_1D of inst : label is "DB9BB7F5E5DEEFF76C0C908380C928C015555400007FFFFE00000058DCBCF0E1";
    attribute INIT_1E of inst : label is "8CCF19DE3BB10EEEEEEEFBB5AF00CC63B1B365833B496635C8D2CC3070EF6F36";
    attribute INIT_1F of inst : label is "47668ECD1DDA33B46668CED199A3B3C6778CEF1D9E3B3C7778EEF1D9E333C677";
    attribute INIT_20 of inst : label is "F615406129B6DB5064A27378D2939B54A0A0A2CAB0C28B25866668CCD1DDA3BB";
    attribute INIT_21 of inst : label is "2A9AC5182B10A22069A01B630B18554E18420421028EED2EECC2B4EAD6D3460A";
    attribute INIT_22 of inst : label is "B4EECEECA5EDF62ECDC473B9A1058FA3854A52A6A8AA86A98AA6A98A829554D6";
    attribute INIT_23 of inst : label is "DF0CDB754366D3BA184A850CC9B0E180DB128B309AB567652F256F2562226265";
    attribute INIT_24 of inst : label is "E9512A2384F6F9819A3128501A142B6D598BD7821542851ADB5662F5E0854309";
    attribute INIT_25 of inst : label is "960B258034B0E9DEDBD6EDABB4B25ACAEE8B6A5B6095C270F3BD336FE3DB1360";
    attribute INIT_26 of inst : label is "ED3BBB60CED08528500DE6E6DB6E834949069EB6362465D6A06AC960B221582C";
    attribute INIT_27 of inst : label is "845F791D8A8DBE50B5B4DC13740C5A26DD5AB52757BD9B5A89B610927ADAD4EE";
    attribute INIT_28 of inst : label is "B699426572C5808E925A502921346F7542BD353EB0CA87406943EB4A994EACF1";
    attribute INIT_29 of inst : label is "69DC33C00A02080B48104050030B0D368D5A1B43684D09852412490196A027A1";
    attribute INIT_2A of inst : label is "1A700428480A13D819D8D60B5050D4057100B17DB6DD9F4EADA3405B9DB9AAB8";
    attribute INIT_2B of inst : label is "2B31D3263A6CE74C9CE9B31D3263A6CE74C9CE9B319CCE663399CCC725263296";
    attribute INIT_2C of inst : label is "CD7011ECC8B062C18B062C14583160C583160C20200001DBBBD0DA34F5D064EA";
    attribute INIT_2D of inst : label is "0532700489D9D6969E31D8482B9453000008E41147218866001326C36C451629";
    attribute INIT_2E of inst : label is "06677604CCEEE1734811559A49BEE9F2D76ACDCB8CDBB6DAE11DBC6B333B9366";
    attribute INIT_2F of inst : label is "766746BEE38596C7566D6E1333B384CCEEE106676604CCECE106677604CCECE1";
    attribute INIT_30 of inst : label is "100000007EC67389FB985876AF0098E1D33810C38F0E8E9E9E9E897303320636";
    attribute INIT_31 of inst : label is "1D7E598F38924832678BC0C0C808B64B7BE58658658658658605EC014497301F";
    attribute INIT_32 of inst : label is "719171B0DAAE62ADCC35311996E623273541C6AA38EDE71CC4FB5D82C7D1C2A5";
    attribute INIT_33 of inst : label is "22E1371C7306ED0CF9F1EE45DE8E398363BB9967B38E60D8EEE47B71C7313CD7";
    attribute INIT_34 of inst : label is "DB4C1C0602472FEF465DC8CFBF1C7313C709B361EE3235C63D1A05DEE338D8E3";
    attribute INIT_35 of inst : label is "D7F499736D960664748ADB6DA3B0C1D5EC065C2E3EFBFAF70935BE4C3316718C";
    attribute INIT_36 of inst : label is "BB5BBDFC819A098F93B87C9976CED27DF13F8387F4FE37DEF66F708837979927";
    attribute INIT_37 of inst : label is "996F48ACFA75040AC160A1011070F6EDDDAF7294146E4FEFA58FF7C6CEFBE367";
    attribute INIT_38 of inst : label is "52E6A5CF6FDCDCB5A633F9B96B4C60C18D89DAD7EF922FEF27AD2977B093BB33";
    attribute INIT_39 of inst : label is "C30C025E986092F0C30097A61824BDDFDFBB7DD6AFAD5D5ABBD65EEB97FCA973";
    attribute INIT_3A of inst : label is "C610E174756F6FEAEB76AA114A4D99B486D832C025C996092E0CB0097A65824B";
    attribute INIT_3B of inst : label is "8B33F96B39DB73DC01B6D96EAA17E69420A7F711BA8A0BB3D75BFCE7FDF9AEAD";
    attribute INIT_3C of inst : label is "36C97B31D4089B270E78A739CE4CB396690442400468AA4667979C1C19193523";
    attribute INIT_3D of inst : label is "11880118852261084210086389210C630804214088C4210021892EC7463C7EC0";
    attribute INIT_3E of inst : label is "84210C2004898C6318C4218E260210086310012261008610000218E248001080";
    attribute INIT_3F of inst : label is "AF3C9A91526A4549A91526A4549A9152624C12644124C8832620C667010C2010";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "0B5A810A4900B492010820154CA480F0F016488D92B38BD0080000059C5E8043";
    attribute INIT_01 of inst : label is "299A1299A1299A1291A12919909485A42521290B485A42421290B485A4252161";
    attribute INIT_02 of inst : label is "7A324D3AF4D9AFF2311092D5A1291A1291A1291A1291D562A8AA288A221299A1";
    attribute INIT_03 of inst : label is "2D755CA3CD1A6699449F09E804E84CE84CEA04EA04C403E00810083DC1B33E44";
    attribute INIT_04 of inst : label is "92F502701A93C067427A01D00E804EA0544944924F48B6F804E84CE8075020B6";
    attribute INIT_05 of inst : label is "2421210908480A8A428A2827149498D4CD964925B6DB2CB2CB2CB2C92CB6CB24";
    attribute INIT_06 of inst : label is "11A285162416CB2CC0110CB4314A16842D2C84A59094AD0B08581090B2121484";
    attribute INIT_07 of inst : label is "290CC4C24D2A78A085802129090848D082621989849A5488842529490849FC26";
    attribute INIT_08 of inst : label is "6D8928B2EAA2CBAA00110532EB265D662349003B4ED8853B7E13E135BE138931";
    attribute INIT_09 of inst : label is "8A4A121292100EAC22029F5A443AB63342225541425085A4D485A4252E81B640";
    attribute INIT_0A of inst : label is "586A9550AA154AA8552DBB76EDC993264C993264DBB76EDDBB76ED92B993E901";
    attribute INIT_0B of inst : label is "2088664622252629A4C21A44E4C9C41880A6030A50C1A911C1450B0D82C161B0";
    attribute INIT_0C of inst : label is "0000000228A24A291452CA2A74E44CD97B3FC858086A33E31326E64CA0908084";
    attribute INIT_0D of inst : label is "0E054D536B6B1225404895012809404A8095012024141506A8A1C90000000000";
    attribute INIT_0E of inst : label is "EDB5C04C2C9A6DB5B6BA13D61A6484D427C132B5641A6AA01A5352710AD6103D";
    attribute INIT_0F of inst : label is "49249249249249AA92097775D69C36C001A514D269B6D72890699204834D06DC";
    attribute INIT_10 of inst : label is "082E8CFAB4D8CC7D098FA136339EF5B104B004924A0220000022220000AA2C12";
    attribute INIT_11 of inst : label is "00315862B18B8EE626378AABD010CD068484250432292B559266993B760EDDB1";
    attribute INIT_12 of inst : label is "109084842421210B421298874CBCCE141D304DE138A29BC2718D4438807C0102";
    attribute INIT_13 of inst : label is "A08208208208208321C2684A6DB9284842C216909484A42521621C0494E30F09";
    attribute INIT_14 of inst : label is "B8AC76AB85CFF6B8AD76AB85830890A4C30A3AF0D5A6D2EE1C69AB1362C006C5";
    attribute INIT_15 of inst : label is "1557A0545149A51485932136C8A1678A29260423D023D020666C5A00211FAC36";
    attribute INIT_16 of inst : label is "2D3999423A51693498CC252CCA520DF3341BCCC01B8C700062B0C563175CC4CF";
    attribute INIT_17 of inst : label is "C5A1C5A98E6CE40812CA14081025862810204B0C1820409650303038892D4449";
    attribute INIT_18 of inst : label is "3140C20008A061000C5030800228184003140C20008A061000473227C9279DE1";
    attribute INIT_19 of inst : label is "A283083A0C5617588208A0396954801A754D3AA6850300004503080062818400";
    attribute INIT_1A of inst : label is "000000000000000000001000045626A24A490984D45449715B48149F890912A6";
    attribute INIT_1B of inst : label is "00001F7FFFE00000080810102020000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "4000000000810008100081000810008100081000810008100081000810000000";
    attribute INIT_1D of inst : label is "5E09B6AD858464236465B19305DA36D0000000000000000000000074D0B04AC0";
    attribute INIT_1E of inst : label is "8A8915122A2EA505050501452804884200205A52A2C190927A43212C94A42C16";
    attribute INIT_1F of inst : label is "C5558A8B15562AAC5458A8B15162A245548AA915122AA45548A8915522AA4544";
    attribute INIT_20 of inst : label is "7F297AE56DA69A64664321267176BF7CA5B4C6DA48531B76625558AAB15162AA";
    attribute INIT_21 of inst : label is "5AF6DA14DB685B7831A38AC91E49DB6F8EC5A766D72A8A2488A14DECF7238536";
    attribute INIT_22 of inst : label is "976A76AF666DB4A8888B39DDE68807C010202698C99698C896BCC9B6BDB2D332";
    attribute INIT_23 of inst : label is "92CE5FFD5176F7EA9CC58B365AB6596859B79BB59A956D3565352D757A7A3A65";
    attribute INIT_24 of inst : label is "B672CE6230C4D965142C10249C09D14A712A560493810264529C4A958125F48A";
    attribute INIT_25 of inst : label is "E472190EECC84A909A94692A28B664F475118C8253210C4338A8224D59922272";
    attribute INIT_26 of inst : label is "4D222252A2A0A20A20204F44924408CCCB259314A466459593448E4721D990C8";
    attribute INIT_27 of inst : label is "455ADA114D0928A028A894A256C816488A142C1189191216D122B02556568844";
    attribute INIT_28 of inst : label is "28E1805183A460070C7661D9D9459A5420474F47A88845663026FA81118AC739";
    attribute INIT_29 of inst : label is "5294A286CECEC6CC8E66266626CECDEF0A140280500A014E38E18E39CF466DC0";
    attribute INIT_2A of inst : label is "12AD8863125AD45E1E50848374F4F1033B0CA099B6D952558DEB5075D9D14421";
    attribute INIT_2B of inst : label is "DA31B0263604C6C198D8339B0273604E6C19CD833198CC673399CCE6BB263919";
    attribute INIT_2C of inst : label is "FDB4F66CE4C991224C9912266CD8B166CD8B176090482C9D12B072BCA6B674E6";
    attribute INIT_2D of inst : label is "81F6B4C38B5BFAFA6C35B0906D24D302417A2592D16DB2FEEA796AD966DD36E9";
    attribute INIT_2E of inst : label is "C7666784888A90DBD936A116912241B0C55A9D2BE893A49771893F6A22D5A4A5";
    attribute INIT_2F of inst : label is "444526A4726CBADFDDF72723B33B44888A90C6666784A88890C7666784888A90";
    attribute INIT_30 of inst : label is "166966E6688445EB7B9CE044CD5090CB9F1A6DB7264C9C8C9E9E9B611A191364";
    attribute INIT_31 of inst : label is "17FFA5EB78190C93250B46C6D8D8B2596BC30C71C30C71C30C666E1B2CB7B05E";
    attribute INIT_32 of inst : label is "591B591A92BAC668EE25633DC4AC6FA5954D64A9A9D40596855A1D4403E00810";
    attribute INIT_33 of inst : label is "36A7D0165A054A4850B0EA6C880B2D02A13AD3B202CB40A84EB6B10165A15487";
    attribute INIT_34 of inst : label is "92687C328E558B2B0F1141B990165A154A491230EB2325172591511B722C90B2";
    attribute INIT_35 of inst : label is "844491B6A5160A22F40492496A2EDBD6E845136A76A399EFDC31360922345908";
    attribute INIT_36 of inst : label is "14929C54C3B0928A9112A898149D8497A515050D20C426CAA20A300D92828904";
    attribute INIT_37 of inst : label is "C9CA804A92AD2C6542A346667AF02492999CE79472E696AA95DE554AE72AAD76";
    attribute INIT_38 of inst : label is "92E62DDCEF9E68E24499ACD1C48935CB894CA4D4EAD202454905FFF559222A22";
    attribute INIT_39 of inst : label is "C21C235C11E11AF4870CD7247866B999C7233996EE25CC5BBCD7477FD1DE8B77";
    attribute INIT_3A of inst : label is "5400604D5B4D4EE6A314BFDE1345C9BDA6DC21C235C11E11AF4870CD7247866B";
    attribute INIT_3B of inst : label is "9A22914DB999529C0D24916C8FD47E94A4955733FA8609A284D22CE4DCA92B68";
    attribute INIT_3C of inst : label is "249272A5D2CC12052B58F5AD6A94A2944925C00835F2BB04559594545050270A";
    attribute INIT_3D of inst : label is "00000118C61B2100002184211D918C200000108E88C61000211D8A974CA852E3";
    attribute INIT_3E of inst : label is "80108421086C8C400086108476C4218C6318C63B610000008C4218C36C200042";
    attribute INIT_3F of inst : label is "A53E01C0384708E01C0384708E01C0384F019670096DE1178070984390846318";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "82CCA4633CCE66799C6799C13A161713403303E4C1986C612100000CC363091E";
    attribute INIT_01 of inst : label is "58F3058F3058F3058F3058F3182CC06603301982CC1660A305980CC066033051";
    attribute INIT_02 of inst : label is "5A7D65DB365A4754C162C8473058F3058F3058F3058F01D84611846103058F30";
    attribute INIT_03 of inst : label is "878AAE30E5A572D472265220DB20DB20DB229332933BFC1FF7EFDB5FD83BEA88";
    attribute INIT_04 of inst : label is "4891499100C844190488244122093309224E24DBD1116D88C320DB20D986C61F";
    attribute INIT_05 of inst : label is "03301980CC0673E31BE3C590C6C6CE431B6C36D949209241A68B6D96D3092412";
    attribute INIT_06 of inst : label is "AC7863C399E926D20B3C3860DC6305860B08C161182C31808C04180823010636";
    attribute INIT_07 of inst : label is "CCF2321911830F16C141B059828C14124B3864E43233063F360B4C2C63B49949";
    attribute INIT_08 of inst : label is "10E4BE4036D900D96F7C79C0379806D3867664C4310E78E6C636636A4624149C";
    attribute INIT_09 of inst : label is "E1630119D9DB783B8BF86061F0C0C3946311166C6030C16316C1460B38EC433B";
    attribute INIT_0A of inst : label is "31DEFFDFFBFF77EEFDFF6EDDBB76EDDBB76EDDBB64C993264C9932447C48FF2C";
    attribute INIT_0B of inst : label is "9BE7333018919086113861131222706E1E1058230E0C0C3C35F2E63B1D8EC663";
    attribute INIT_0C of inst : label is "0000000B8E1B238DC708E38D26973FFC3ACB4C1663A06838C8903122124E1E73";
    attribute INIT_0D of inst : label is "01BABAAE8E8EC196AF065ABC15E0AF055E0ABC1782C015715634C9A000000000";
    attribute INIT_0E of inst : label is "0DB666B1B2F3CDB1B6CC6C18F3C6641C3D8348C186F3CE009D6875C947B7F307";
    attribute INIT_0F of inst : label is "79E79E79E79E7A555B2F33370684B6D000BEDA9BCF36D9B8C9CF19264E79B6DC";
    attribute INIT_10 of inst : label is "E4B16E43CD2E10C61B18C3638104A65CF3F6364925B9BB9BB9B9B99B9BB518DE";
    attribute INIT_11 of inst : label is "FA9C9D393C64B09396C4E557C5824560C0460231D58C82ABCB09A4C48931221C";
    attribute INIT_12 of inst : label is "D82CC1660B305982C3018E39D8C2C28263617B234E78F6468C9400677F83FEFD";
    attribute INIT_13 of inst : label is "38E38E38E38E38E404460C04D3620C1460B3059828C1460A301A64035ABD030E";
    attribute INIT_14 of inst : label is "61999C0E1752AC61999C0E174C66C63D0E7B03919FBC8B9B64EC0E3E399E7C73";
    attribute INIT_15 of inst : label is "CAAF96B5BCA46FCA32489C98261CE1B79491B99CD6DCD6C15BC73364CC3519DC";
    attribute INIT_16 of inst : label is "858D41681D6AC4B2596A45B6AC5E399EEC737BB6FE4FC9B5393A7278C91272C9";
    attribute INIT_17 of inst : label is "0B470B4D963B82C5880B96C58B10172D8B16202E5B162C405CB7E7E86085C320";
    attribute INIT_18 of inst : label is "CE6F496EE737A4B77B9BD25BBDCDE92DDCE6F496EE737A4B773D9BDCF59D7347";
    attribute INIT_19 of inst : label is "E4CF2CD33C9E5A7982A0AA994C36DDDB6AADB556F9BD3B77B9BD25BB9CDE92DD";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFEFFFF89E63716F6D8C81FCECCD83A06D36C56D90DB10";
    attribute INIT_1B of inst : label is "FFFFE080001FFFFFF7F7EFEFDFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "BFFFFFFFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFFFFFFF";
    attribute INIT_1D of inst : label is "2474693E1714F9AFDB181C287221C1B02AAAA83FFFFFFFFFFFFC00C2E3424007";
    attribute INIT_1E of inst : label is "46648C891990055005500158C4F0463124B97D6B11275B49050EB6824A30B0ED";
    attribute INIT_1F of inst : label is "232246448C89191232246448CC9191232246448CC9191232246648C891912332";
    attribute INIT_20 of inst : label is "BAD2CD101B3CF3D3D1BC8C111C99C0C2526A39A1A728E68D3832246448C89191";
    attribute INIT_21 of inst : label is "AD1B25896C93ADCF8F5CB92E697274B8E37AD9B968C645B2444CB6095ACB625B";
    attribute INIT_22 of inst : label is "40E38E3895BB122C4475FEBE1977F83FEFDF9947BE4967BF6943BE4B42C96C5D";
    attribute INIT_23 of inst : label is "DB399E3E5EC8F1E2E372F5CB70E10407B66CF66EF5EBD2839AC3D2838787C79A";
    attribute INIT_24 of inst : label is "F1582B9B079795958B136CD9F3B62D6D158B1C41BD66ED9B5B4562C710EF4B2A";
    attribute INIT_25 of inst : label is "0984C26336922ADAF0C4C48B12E9D959766D7BB96AEDAB7AD6BB9179CD9BDBC4";
    attribute INIT_26 of inst : label is "3811116ACAC81881081B3F62DB7C042B2B82DC57166F7756EDD9389C4E252713";
    attribute INIT_27 of inst : label is "94716488BC45B81D97B2DC0B762EC96CEC89176532688B59C5B00DB6CB5BB222";
    attribute INIT_28 of inst : label is "16B3362D66C89DCC71494C2525952B7ECD9DB5B792D997D9A4C979765B2F9CFD";
    attribute INIT_29 of inst : label is "645AB1397979796B6B8B8B8B89292F364489312626C4D8B8E38C30C736B8B693";
    attribute INIT_2A of inst : label is "DAB2F79CE4EF7B71F15C625E8F8F8D8DAEF2BF08B6D88BD6C5BB98D977D8DDB5";
    attribute INIT_2B of inst : label is "3BE7599CEB339D6673ACCE759DCEB3B9D6773ACEEF77BBDDEEF77BBC24BDE6D2";
    attribute INIT_2C of inst : label is "4C3189BB93A74E9D3264C99BD7AF5EB972E5C886433192DDDACF0AE736D90E35";
    attribute INIT_2D of inst : label is "6F3431BCF4360181A59190D8867FBE998C8CF86D67824D2698CDC386D9B3ED9F";
    attribute INIT_2E of inst : label is "3222226E64464B721CD9C88CDC95CF27962C458E0C5E16DAEB70E4D91131B736";
    attribute INIT_2F of inst : label is "2222DBDB5B92418644E1F67991192E64464B3222326E64464B3222226E44444B";
    attribute INIT_30 of inst : label is "C887887924D62BCB1EF36023B88E47143358C208D1A3E3F3E3F3F41C4DC4C883";
    attribute INIT_31 of inst : label is "C80BD69F86743A489066393136366DA4C69861C71C7186186711B94493487F30";
    attribute INIT_32 of inst : label is "65A565A4D832791633113CC6622798E2DAA1B6543604064965460DBBFC1FF7EF";
    attribute INIT_33 of inst : label is "4AD8101925853A364C8E6CB3680C92C2891B2C5A0324B0A646CB0D0192595183";
    attribute INIT_34 of inst : label is "5B6F178C789645ADF0889E02501925951A33061E6CB0B2E4B25AA9864B12C0CB";
    attribute INIT_35 of inst : label is "E2365ADA35DC66CB1DF85B6DBB11842C1657588F4ECE729725E5E4C6BB0624C4";
    attribute INIT_36 of inst : label is "86DB395C66161B2B7648B26EC6F0B6D930D6C5B1B796BCACCDAECDF041313776";
    attribute INIT_37 of inst : label is "6411C7845EB65393BDDCF898851816DB652B5FC31D96DCA2C3E15171F8A8B0F9";
    attribute INIT_38 of inst : label is "5C78B8F1765B061B610CB60C36C20A142DDDB786312DD9676DC35718E5B11911";
    attribute INIT_39 of inst : label is "6CC61E1B6630F0CB39878659CC3C367396DEF65870B8F171E6E5BCF3677B6C38";
    attribute INIT_3A of inst : label is "67B9BB622F7973DADE576A333E39F63C3986CC61E1B6630F0CB39878659CC3C3";
    attribute INIT_3B of inst : label is "2B192D7A45251B73E0B6DCC11206C421084EEE48C9C9F7BB57DB1296228DE5EF";
    attribute INIT_3C of inst : label is "16DBC99B297A5B978E76A739CEDB3B677FF0FFFF8059EE222256CB5B5C8C9191";
    attribute INIT_3D of inst : label is "210842004230631086310863189080000042108C484000842118E66CA11225B9";
    attribute INIT_3E of inst : label is "00000001084084000840008422C421084218C63061000000084218C224631884";
    attribute INIT_3F of inst : label is "1A92224448C919232464889112224448C9196991869222088811931890800108";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "821880231C4C26389863898528163211C070094403802AC00100000C0156000A";
    attribute INIT_01 of inst : label is "4851048510485104851048510824412209104880440220910088044022011048";
    attribute INIT_02 of inst : label is "7275759B365A472151264045104851048510485104856158C6318C6301048510";
    attribute INIT_03 of inst : label is "424AA93C91E548C2496E09600160496001620162010000000000137998A2640C";
    attribute INIT_04 of inst : label is "013100B010A1C04B001800C00600160032E72E4B4B0B24B8496049604B025C17";
    attribute INIT_05 of inst : label is "08108084042023510B554743A6A6AD400925124B2494492810580030006000C0";
    attribute INIT_06 of inst : label is "FAF466A149A490005B3AEA238A21040208084101082028824410082021040572";
    attribute INIT_07 of inst : label is "44E969149142841E412B9040820410124AB452D22922853472080A6A2110B825";
    attribute INIT_08 of inst : label is "28509D204A748129ED6A68A04BB409714E52A4A228856BAA5C12C1212C129C8A";
    attribute INIT_09 of inst : label is "D121008B4B4FE82B59745050E8A0A1552111322C2000410112410208126CA11B";
    attribute INIT_0A of inst : label is "1142C4588B11622C45A922448912244891224489122448912244892C7221FF7A";
    attribute INIT_0B of inst : label is "89C631291541484503105031211720E41C087122854A0A281DA0522110884422";
    attribute INIT_0C of inst : label is "00000009451A9144A28891448692AFF82A53440221200111A44A289112450E73";
    attribute INIT_0D of inst : label is "0192A8AA4A4AA952A6A54A9A94D4A6A54D4A9A9352554029552A818000000000";
    attribute INIT_0E of inst : label is "049572A8AA51449092AD2A14D152E40C1F8328A142D146021868354146A51101";
    attribute INIT_0F of inst : label is "20820820820821554A67333506849255559C5A094512559A5B454B72DA28B24C";
    attribute INIT_10 of inst : label is "C4B16D43A485485C090B81214041090AAAB2044927DDFFFDDDFFDFDFFDB50AC8";
    attribute INIT_11 of inst : label is "025A94B52AD49009444051574586CD2040020810910A02ABAAA494A24528910A";
    attribute INIT_12 of inst : label is "C8004002001000820100051348C28242612129612D5452C25A94002000000000";
    attribute INIT_13 of inst : label is "14514514514514520DC20400492904022001000804402201100A200A1A1F060C";
    attribute INIT_14 of inst : label is "2108840A1540042109840A1544364D349A3342B09F340A8B20CC0A2A149AD429";
    attribute INIT_15 of inst : label is "A2AE95ACAAD2ABA96A255A48510AE1955A4A9095801580014942932C4C200884";
    attribute INIT_16 of inst : label is "8C930B20B86A4592C9986CB98ECE7932ACF2CAB67A0F41ACB5296A55A9012880";
    attribute INIT_17 of inst : label is "0C050C0D1D2AA2C5885932C58B10B2658B162164CB162C42C997A7A8608CC320";
    attribute INIT_18 of inst : label is "A8245864D4122C326209161931048B0C988245864C4122C326358A15C1155105";
    attribute INIT_19 of inst : label is "6C656641958AC82BA800AAB04D2249C92AA4955260917326A09161935048B0C9";
    attribute INIT_1A of inst : label is "000000000000000000000000018AE23127248581FDC5C4870125724064B0C912";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0450213C151CA1ED032008707000A2881555540000000000000000C2A3424040";
    attribute INIT_1E of inst : label is "46648CC9199005555000015CE5A846316D9B3869912549A5468A93494D38E0A4";
    attribute INIT_1F of inst : label is "232246448C89191232246448C89191233246648CC9199233246648CC91992332";
    attribute INIT_20 of inst : label is "18124E0009145111423A081208888044002C308022B0C2111432246448C89191";
    attribute INIT_21 of inst : label is "2C1A058B68162D0D4D5AB1640B2045A05322E19130C645A04458940BCEDA62DA";
    attribute INIT_22 of inst : label is "09A61A61B5A912244445A8943100000000005B06B40B02B40B02B40B02816050";
    attribute INIT_23 of inst : label is "496A1D2A5050E14281224489C1828A22008C428C41830011001100110D0D0D00";
    attribute INIT_24 of inst : label is "73586B490692B0B48B126ED943B76D25148914C33176EDCB49452245304C492A";
    attribute INIT_25 of inst : label is "0B0582C3B6922A4A5045C48912A95B59524E7BB12AECAB2A529B9128C7091946";
    attribute INIT_26 of inst : label is "2811112A4A58018098823522493C226B6A424C7313463552649960B058252C16";
    attribute INIT_27 of inst : label is "B4516C8CBC449819979248092664CB264489126DB3688949C494099249CB3222";
    attribute INIT_28 of inst : label is "129A362534CDC99C414948256515293ACD9494971655B38CA6C971264A2714B8";
    attribute INIT_29 of inst : label is "244A91636363636B6B1B1B1B1B6B693C4489B13626C4D8B8820820873C01931B";
    attribute INIT_2A of inst : label is "5A92D6B5ADA52B51514C621A9A1A0C81A8EA9C4C92488972C4B908114548DD95";
    attribute INIT_2B of inst : label is "39AD5815AB02B56056AC0AD5815AB02B56056AC0AD56AB55AAD56AB424B5A252";
    attribute INIT_2C of inst : label is "48640DAABA3468D1A3468D1B162C58B162C5890D0683425CCA4A8AA71E59284C";
    attribute INIT_2D of inst : label is "CF246430408080002591804806FA28B41A0DE0816F040E24BA07060802328194";
    attribute INIT_2E of inst : label is "632232CC444443221211CC8C4C95CD6293264C8A244A924AC230A55911331222";
    attribute INIT_2F of inst : label is "3222C95B5123650ECCC3FC7111190C444443622232CC644443632232CC644443";
    attribute INIT_30 of inst : label is "C44344500452214A32D16022AAC4261872720410E9D343434141401AC5AC4513";
    attribute INIT_31 of inst : label is "2209869F0E5229254A62B4B28644000052B4D30C30C30C30C721ABC840012E94";
    attribute INIT_32 of inst : label is "24A524A648321086131108526221024262A4B354970402496404848000000000";
    attribute INIT_33 of inst : label is "4A4C1009258030170E1A259B280492C01C0966CA0124B0030259C50092590121";
    attribute INIT_34 of inst : label is "49E7279020D245A5A0889452D009259030164C8A24909064904AAC8649124849";
    attribute INIT_35 of inst : label is "73344ADE7CD4D6CA09E24924B9128865361249055A5EF7BC45A4AC47999224C4";
    attribute INIT_36 of inst : label is "42497B4C6206096976489664E250324B10F2C4E8969295846CA6C9E081B1B672";
    attribute INIT_37 of inst : label is "30B9C6044B966343B1D8F4544E0892492F79CF03209C48C301436180A1B0C050";
    attribute INIT_38 of inst : label is "D021A041C271A45923061348B2461C3864911283392D993224C1469CE4919911";
    attribute INIT_39 of inst : label is "7D820A13EC10509F608284FB041422529C4A525020A04140838DB5A6656B6810";
    attribute INIT_3A of inst : label is "73BDB3322D2933DA4E5320173A21C438A083D820A11EC10508F6082847B04142";
    attribute INIT_3B of inst : label is "39192D2A4D2D1133D492484310028A73182CCCC4889DA699534996932688E5A5";
    attribute INIT_3C of inst : label is "1249491D202A499244268210844B91723FF07FFF9048A22232724B4B4CCC9399";
    attribute INIT_3D of inst : label is "0000000000010008421084000000000000000000000210840000E474839726A5";
    attribute INIT_3E of inst : label is "842108421085086318C6310840000000000000000218C6318421000420000000";
    attribute INIT_3F of inst : label is "021614C2981302604C0981302604C098130200303000606181B0A10CA1084210";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
