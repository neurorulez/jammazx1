-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "066F2D985C0060208D0013EC8455004240028FB3723A3CFA7555DF4B75E7AE55";
    attribute INIT_01 of inst : label is "67845B67B19FB6664B71A2B65AEF917578099D2496965D279F4898BF0F400030";
    attribute INIT_02 of inst : label is "8923BCB734C2C42F7BEC0F178006879B03D8B5E216F800000016A39022AB7C8E";
    attribute INIT_03 of inst : label is "ADD0BA773FF9B098F788D179FFA929F20DA4135ECBD9BDCD9CE63EDB7DB6766F";
    attribute INIT_04 of inst : label is "6629CA4825F10EC3476320998924E484FDA18B622BEA468EC6A747B1A9BFFEDF";
    attribute INIT_05 of inst : label is "F3594EC40006E80008FD00382CFE20D928718C8A111102D2A6A53283437D3AFE";
    attribute INIT_06 of inst : label is "E79CF3CF3B73A19023C8783E4F91FF832C16E6F33A7CB366285C4791020A3273";
    attribute INIT_07 of inst : label is "B08A15800B0C97E57547EABAA1A4DE201323A97A96283F9801948E919288197C";
    attribute INIT_08 of inst : label is "000818D38EA344A51A462C9F76DB249362144FE80F7E108C52D7380C525BC924";
    attribute INIT_09 of inst : label is "46DFF6E3AE597E4E32E6EFAF4DA8C6C6DFEBE6A111FE8CA18812FCFAC05979E4";
    attribute INIT_0A of inst : label is "F0CCE11568836291A1743B11F99B6DF02002407DCC0DCBAAAAD25FFDA2D77B41";
    attribute INIT_0B of inst : label is "2205FEC24CFEA6E1E2504D893DBBFDBF9C720A00319419FBF7FDEDCD3340C299";
    attribute INIT_0C of inst : label is "8022319B1454888993C8FB6206DCF1366A004881502115ED17BDA00DBFF65B6D";
    attribute INIT_0D of inst : label is "7E91240278318886A8294D8A42A94837EA69519B42E4FE2913DAF91628A50A52";
    attribute INIT_0E of inst : label is "9DA062AB23DBD0AC359FBE3FEAA67DA03CA73749F18BEF18660F9DF33F61F7E0";
    attribute INIT_0F of inst : label is "B9187C3323F6922A04233D63D647D867D2767B1EB23EC33E93F2C0FB0FD619F4";
    attribute INIT_10 of inst : label is "01AD77F0E4000B4B555D76EBB75DA0844ADC9C90540845B929911FB591540845";
    attribute INIT_11 of inst : label is "A0644AA819127BEE05FB7F4BCBC82540B93FA6FF9BA71A14F41808B2024B198B";
    attribute INIT_12 of inst : label is "4632C57DBD8F05F1624E00D2BFCB013ABD130F221984D81CC26C0E7200A9B1E2";
    attribute INIT_13 of inst : label is "08020AB9CEB3D5E2B12F17D79F446782110885086384899E4D15691EB29D8971";
    attribute INIT_14 of inst : label is "F82345B7061798208049ED26FC0104021842A000936708B91D9810424400082B";
    attribute INIT_15 of inst : label is "B8084F8272109F00E0023E09C81D9450007CA2C013E514011F28B10CF96BE219";
    attribute INIT_16 of inst : label is "96937B1B00410082436892A66830012EF24716D992AB3A9090D1000805A54777";
    attribute INIT_17 of inst : label is "16C43600130082AEAF4EE61CE45C33E4626D62636E94D8D76D04A0324492D6EC";
    attribute INIT_18 of inst : label is "AC6934A8814A8DC7D2947909BBE5DD84F452147204868875350C08450A2BEEFA";
    attribute INIT_19 of inst : label is "229A48F9B9FBECAAA480606D86BD4D81489B0C1122411DAEC76BB1DAFC7F96A7";
    attribute INIT_1A of inst : label is "AEDD8B79E284932BA71C9172E8370FCD0654D4202080424C9CB8E9238E922A69";
    attribute INIT_1B of inst : label is "DCE4C5DB0D83E29E49D908214BAFFCC1FFFFFC3FFFFF0C01999E05E9934E9F9D";
    attribute INIT_1C of inst : label is "F3CC9FBE3ECA63AE1219ECC3EC2377E1390CFE0F32B306C8048AD46B6DC924EE";
    attribute INIT_1D of inst : label is "B9249D7E8CA0C40D5210254D59071345934764C46C9256A88975184BCA052063";
    attribute INIT_1E of inst : label is "83C050259CC6C9C632002B37C1A4E9FBC001479157427BC930F4BF5F114F9D6D";
    attribute INIT_1F of inst : label is "9D3E637893A97AF8DF8E7F6494336A44838871344B0A34003FA2ADFFCC1E70AD";
    attribute INIT_20 of inst : label is "FD5FB396C4F9E56352E6CF2BB84C4194BEE674C19C48704D58E89AB1D1063A62";
    attribute INIT_21 of inst : label is "803FFFC7803FFFF87FFFFFF87FFFC7803FFFC7803FFFF87FFFFFF87FD2AFFBAA";
    attribute INIT_22 of inst : label is "B54AB54AB54AB54AB54AB54AB5457F32AA97872C500DA403C3D3D07071E9E847";
    attribute INIT_23 of inst : label is "09290600208087AB5555AA55552AD52AD52AD51AB54AB54AB54AB54AB54AB54A";
    attribute INIT_24 of inst : label is "8B624831F02480093701009D40DBC7C0BE9F87E05FBF0E2600A849B60118C80A";
    attribute INIT_25 of inst : label is "D00640015158D55428BA00DDD6DFFEF400082384DC4404084601801044600411";
    attribute INIT_26 of inst : label is "A007E0BE73649954C921D9083A27A8B5B6D121D7E859893B5D7483B250CC392B";
    attribute INIT_27 of inst : label is "A555AD9C00ED258FE3496E00736B554AA555AD9C00ED258FE3496E00736B554A";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "D10A5CACA0E300C3E538897D8E8E09D5001990154A1F68588FFE7F223E63A773";
    attribute INIT_01 of inst : label is "E80692480A21D7C07A78844736DFDD179D5BA59DAB65324028958D00A200CD80";
    attribute INIT_02 of inst : label is "24A75EFFB5A340F9468F5ADCA00213AC7371FEE43F990000000D60166E392282";
    attribute INIT_03 of inst : label is "B799D33092FD280567520471E67A8858DEBDB57F981EC9E050F0490411607C31";
    attribute INIT_04 of inst : label is "027A49E0F1F317D1A7AA72AAA8700DFB8115908570214ADCF29B6A3CA2849386";
    attribute INIT_05 of inst : label is "F638AFAA2FAA5BFBF7117F527FBE62FA3A7C7E5BDA081724484952F1BD528EA1";
    attribute INIT_06 of inst : label is "48A91490125172A019AF8A4290A20077FDF1B0BF7BF5DDCB4ADD57AA9F1D7639";
    attribute INIT_07 of inst : label is "91D178C9524001C9799DECBCCC82679657F8CF63362DC0CC6F3A7DDE01E88A05";
    attribute INIT_08 of inst : label is "E5B1F1A4E03D10BDE885EF377965CB2042C3B88AB2004ED5571D5E5550E21B41";
    attribute INIT_09 of inst : label is "9500090748A00090748D020090000381D4924B6A324BCCC655A20252AAEAAB4B";
    attribute INIT_0A of inst : label is "E29D04E247151FC2BEA35DDD0AC4184BDB7FBFE95454503AC36FA4A8450A908A";
    attribute INIT_0B of inst : label is "444000D491632EEAB41952840929492E46B55C5F44FA30C1B32E494A4464A92B";
    attribute INIT_0C of inst : label is "FE399A46A2AE5270401600DF6836025390F2A54EB95DE2422948450A0006A488";
    attribute INIT_0D of inst : label is "F12A136C014B0E733407247F1AD7A9502000222420090875AC231937FDCC74AF";
    attribute INIT_0E of inst : label is "441284C25C92DF41820C1BE43F4A891B4BD5CBA2293254A398556148884B8374";
    attribute INIT_0F of inst : label is "6C5280CD54A108572BBC485524897685451092A9244BB42A2884A92ED124A151";
    attribute INIT_10 of inst : label is "18FEA1750D9655BDDE92489244927F6DBE362143AE57786C4662250846AE5778";
    attribute INIT_11 of inst : label is "72B28F5DACA6924A50048452B0116A2802422A5214A9C37156108A3FFC99C194";
    attribute INIT_12 of inst : label is "150295EFB4EAAACCCE2C598875D52A8EB9B6AA4A8AD92D8525B24006B3E2CB0D";
    attribute INIT_13 of inst : label is "C8084370A570F3B9735AEEEEF8C9EBA28160B38B21A01A3C05462038F35F57F3";
    attribute INIT_14 of inst : label is "1A35D3635CD9D7967A26C0136EB6DB7FF70EE14E4821A50FB40E4FB7AC00090F";
    attribute INIT_15 of inst : label is "7B0800D5D60081ABA820035F5611B9D8020DCFC200EE74008373E0003BC7C000";
    attribute INIT_16 of inst : label is "6009B076ADB6DFFB27E800EFA0AAA88DC64B16E4EB573D7F6B2B6FB6AC33BE13";
    attribute INIT_17 of inst : label is "818507C6815B6AA2A2FF9F9EFACB71851E8C1E54450E031C358CA00067419886";
    attribute INIT_18 of inst : label is "1B00007D4EBDA1D12FB4D40E284D00830DAFED45EB595A151507B6A3DDC2C262";
    attribute INIT_19 of inst : label is "389B8E11111249AA0925AD32DEFC92D8E66C9B0990A8EB552A9D4EB542A52DB5";
    attribute INIT_1A of inst : label is "399E7CD7A1E02773ECB656752B6B746167D45416DB6FFFD99EE8DE388DE38A6E";
    attribute INIT_1B of inst : label is "557433AE2F1FEF15547EE5A5F41000FFFFFC003FFFFCFC0181FCE70840800013";
    attribute INIT_1C of inst : label is "849D0C1B739EFC02F7ABED54BB4404E557697BA12AD2A44894881A2CB2B2C820";
    attribute INIT_1D of inst : label is "5659040BCCC64164695399D311D1BE7394D3078D1A4926CD11EFD9753B27A228";
    attribute INIT_1E of inst : label is "B18B1A91F5FDDEF56B6D35454A8A30C196BB2E37817EFB5F4A25BC44B8956596";
    attribute INIT_1F of inst : label is "3DFEFD53A8CB78A50400B101BA247BE6D1A14812AD03900005D6D120199C0108";
    attribute INIT_20 of inst : label is "D73FD99A102E428456B7FF5FA950D7DF288090C8D0DD4469DEF253BDE727BE42";
    attribute INIT_21 of inst : label is "AABFFFD2AABFFFD52ABFFFD52ABFD2AABFFFD2AABFFFD52ABFFFD52A9772AE7F";
    attribute INIT_22 of inst : label is "2C66D3992C66D3992C66D3992C655B1FFFD524E4CDB4C6A9571F1D5AD58F8F52";
    attribute INIT_23 of inst : label is "40820200208085C66C9CC9631B4E64B19B4E64992C66D3992C66D3992C66D399";
    attribute INIT_24 of inst : label is "80000100F9000D5CE111940DFBD41FA0BE5F99E25F3F333649C6335E7A0BC44C";
    attribute INIT_25 of inst : label is "12C8DAD4A2ED29BDAA9C03CA39325A88012101E035240564A64992420A649083";
    attribute INIT_26 of inst : label is "200700053380A52135B8116EE05519FA879A6A08CDA358A8D3FB0073D8B86535";
    attribute INIT_27 of inst : label is "633364B55549B9F01F3B25555A4D998CC666C92955A49C7FFC724B552926CCC6";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "5025B83738EA377DC33A810832B576F400108F00254BF20ACBAA2D334A410201";
    attribute INIT_01 of inst : label is "EC369B7B1B3744090C4000062A8FDE07D7FBB99DB4D64B2EDACA320AA22F7507";
    attribute INIT_02 of inst : label is "36A77E7FB58E5C94824A229A4000A6AA3C43F8E2FF180000000A34346E209152";
    attribute INIT_03 of inst : label is "4672CE42003B8404C3540602E5FA925AB5B5637ED41031090284045146B4540B";
    attribute INIT_04 of inst : label is "2070C90081F00081152E72BAB8700D8043A14341443A4392E76FC939DB632C48";
    attribute INIT_05 of inst : label is "F6592A822ACFD0952A19527AFE3E001130552E8A90D198B66E6D70A1092D1E5E";
    attribute INIT_06 of inst : label is "6BAF74DB9B718BB391A53A6E9BA3B02F8856302A7FFA3D0F6AFDDBB0B7BE2BD0";
    attribute INIT_07 of inst : label is "E65694FF506001C1AE0110FF00A007144384F023C346819C12B4AE94862D8A5D";
    attribute INIT_08 of inst : label is "C5B95587C6A1D2D96E9649A03FB7FDB1578804CAE3846085FF1F7C75F0E01BC7";
    attribute INIT_09 of inst : label is "C5B60DC772B360DC772D9B6CD8618282A6DB6E85027542611DBDDA282AC2830F";
    attribute INIT_0A of inst : label is "E3DDC6037896CA2734E750661B5A61A0A000096D9E5B19B9E6C826EF658EDECA";
    attribute INIT_0B of inst : label is "666D84D6DB93AFEBF61B58D00DB0ADB98EFC0A0167112366EE736DE3676245BB";
    attribute INIT_0C of inst : label is "A6D31B5833B45AA4609AD3092CC73BA79C56F85AD369437B2D6F65AB6C26B6CF";
    attribute INIT_0D of inst : label is "A5BE074FB961B4E395CF03289CC02876A800333776CD8C60B5353FC2A36FA6C0";
    attribute INIT_0E of inst : label is "8C32D6DB68DB8A4182366EA9FA6CCD936F87CF033DB27433EA5AACAB1C74CDE8";
    attribute INIT_0F of inst : label is "8EDAD8F476E99E5A6D286F69B6EDC6D2C630DB4DB76E36963186D5B8D9B6B4B1";
    attribute INIT_10 of inst : label is "385C01F58D145652CC1A60D34698000502C76CF6B4DA518EC7ABB70DF6B4DA51";
    attribute INIT_11 of inst : label is "82F40D60B5069B6E5B66C65A90196B6DB3632A2B766F8A0EBEBA200001B9C035";
    attribute INIT_12 of inst : label is "6EAA188F25C55479CF6C519CC7D72B1FE117BB4F8AFBE68D35F7C406A20A8125";
    attribute INIT_13 of inst : label is "8802004CC2721B9370182E0E10C16D168B45A15E207001010167800030550477";
    attribute INIT_14 of inst : label is "1F9B7CC7D3E1D2C9240D6D0035010010129C794CAABCFFC5F834800034000802";
    attribute INIT_15 of inst : label is "DE31C8AB5C739156BCE422A579F3E013DE8F019EE4F80EE627C036351FB0E429";
    attribute INIT_16 of inst : label is "D680190040400400016D00EEC381E80A2B420A014DB3A00252C3400844811B7D";
    attribute INIT_17 of inst : label is "B6AD041A809087EBE82F4C50C29450D2A588A56C6A40611281F59C58E86E6E8C";
    attribute INIT_18 of inst : label is "1B0801884201A5F680B400E4297D09815C000D7082961EDF1F90082C08CB6FBA";
    attribute INIT_19 of inst : label is "C0F7F01DDD9B6FAF1F7DC61AEEFC1AFDE07DFE5D8090150A850AA542A1552A31";
    attribute INIT_1A of inst : label is "309094562C402AAE29151074C8675945147C7E402002005AD4EE4FC0E4FC1BDF";
    attribute INIT_1B of inst : label is "50F4671E2F17E84A58F8C0A103A00F01FFFC03FFFFFCFC001E1C761C20210481";
    attribute INIT_1C of inst : label is "46DDB66EA79FF16F37BBF5D6E37651B9754DFB2D18F105441C60103FDBFF6C4A";
    attribute INIT_1D of inst : label is "7FED8935426259C44211A3F6B1C19D03372925F83CB3A0639052C52B1308362B";
    attribute INIT_1E of inst : label is "319E90A35F4F70FF8FE737D2CBAC7366F73A2CB437E7FDDF62F5FE45C4DAAFFB";
    attribute INIT_1F of inst : label is "37FFF02CB1EBFCAF9AB2FE43B0BD7D5654C2F004257212AA87C8A4401D0021CE";
    attribute INIT_20 of inst : label is "2DAAB79CB1BC72C74232AF658958049294629A15000D276594A34B2941052B44";
    attribute INIT_21 of inst : label is "403FFFF1BFFFFFF33FFFFFCCC03FCE403FFFF1BFFFFFF33FFFFFCCC010A80080";
    attribute INIT_22 of inst : label is "3C7EEFE7C38110183C7EEFE7C387DBFFFFF9C41C3DB907C295D1D26232E8E8CE";
    attribute INIT_23 of inst : label is "00DE125165C5930183E3F77F1F0E044060F1FB97C38110183C7EEFE7C3811018";
    attribute INIT_24 of inst : label is "3054008810805A7268670C0C93F4206DDA4F0006ED1E031403460308C30B029C";
    attribute INIT_25 of inst : label is "119C218254F1943D1B40000C0FEFE458000800704A0402002401001012400405";
    attribute INIT_26 of inst : label is "1007EDBC794701A1AE6D1A4CC002DFFB16FB6B8D49242A6A51000E241F8B31DB";
    attribute INIT_27 of inst : label is "B5A5B6D9998E3E0000F8E33336DB4B5A52D25B64CC6383FFFF838C664DB49694";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "4825889F18BC277CC6AF411BB11276488030D5E6354AAC7A10A2C8624243C301";
    attribute INIT_01 of inst : label is "05AA492A999568C13E88022E06B7D4B55BB8104C9ED659B5924851EA028F7617";
    attribute INIT_02 of inst : label is "9B04E0775C6D99C08211098060040278304288E4D11900000019B5254E509552";
    attribute INIT_03 of inst : label is "84F19E239B637449CD1A98E7798986B4D729A65F10226A296215805145950B1D";
    attribute INIT_04 of inst : label is "30676D3C960A91B020D50351500D6644FCA61301D7DB0F976D27CBDB49334C4F";
    attribute INIT_05 of inst : label is "F3962143B22C86D5A3F01A4EA2035226A78BA590E3F559972F2E7F10222B1056";
    attribute INIT_06 of inst : label is "AA754D52C93CB91B7025A7298A6120AC9B56A20607796005A220D790B2BA2065";
    attribute INIT_07 of inst : label is "B6220124126B05CE2C08FF3804204A504D11FC5C05223EA8C992B6672A050DD3";
    attribute INIT_08 of inst : label is "E0FCE8C607C67E20D3F58478049724B1B42C4F81E1F83318A0DA2D68A01ACDBC";
    attribute INIT_09 of inst : label is "F993EC8232B93EC82329EF2658B6FF6D4359EC437B36716F0FB9CC2A6059F98F";
    attribute INIT_0A of inst : label is "130D83312BD768EB8467395491586180800009248CDD88EC936ED2657DC64AFC";
    attribute INIT_0B of inst : label is "6364F882DEF98B03A62D9FD00498A49F0866C6CF71C339227C7524F1632C44BC";
    attribute INIT_0C of inst : label is "A4C3015897134ABD008AD3096ED511E4183AC8585B2E712BEF257ED327C416E5";
    attribute INIT_0D of inst : label is "C4B7034F9B71306059C605A3AE2033369DC81116F265F80CB5A820048DA9A2C0";
    attribute INIT_0E of inst : label is "8AE2F2092E49EB3A5C922649712E64AD6492842B9C9A3C99E8DFA8AA112244C6";
    attribute INIT_0F of inst : label is "AA08D5F53249924B65CE2524B2E480E2B628492597240715B1424C901CB238AD";
    attribute INIT_10 of inst : label is "9890F179E55CE6D688D822D1560A820902D5059616CB9DAA2FA9920D9616CB9D";
    attribute INIT_11 of inst : label is "9A74E6279539C9274932FC0E8AC933E4997E042B068C0C4017DFFFC00248D356";
    attribute INIT_12 of inst : label is "1DB42BA17B4532EADBBD6785D1E723114825D5B482B6DB015A4902B36A4B8134";
    attribute INIT_13 of inst : label is "882B60488A3159442A8D0747404C20744A050050B300459800B180A32C428402";
    attribute INIT_14 of inst : label is "07F7B744DE481A09241B7D02314000101AAA1D0F236F730550F6024824000D82";
    attribute INIT_15 of inst : label is "960008294C001052980020A53C026020009300001418001020C0000107F88001";
    attribute INIT_16 of inst : label is "BE811F4D50000402405D00667373E051B21F0A390FA24E024642C04047A50BED";
    attribute INIT_17 of inst : label is "D62810DA00940549490814E7C3F338CC5782568409F44D2616C0E03C1BE7DF09";
    attribute INIT_18 of inst : label is "314A1288D7017F960091A07E13BADF614DC00BA48232176A8A824034086D7DB4";
    attribute INIT_19 of inst : label is "01A8004CCCC925BFE493C66D33BDED26CCDB60EF3080562B1582E170B8584354";
    attribute INIT_1A of inst : label is "D04358260CE012B85F5E07F9F33A6FF078AA2A080002014CA2FBA001BA001EA0";
    attribute INIT_1B of inst : label is "AD886FDA3D52F18A988E47CE2A88000000000000000000000002AF85402A05A0";
    attribute INIT_1C of inst : label is "024D9226470910249B3C1D864273F18123245DDE7167118C58E462824B892C7E";
    attribute INIT_1D of inst : label is "71258FF6716E1AC08A67098A9EA3C8836A21F020BCB7796B599CA2A771701433";
    attribute INIT_1E of inst : label is "D0BE2609450500500F76C7B2AB2C4922731BA0E8921207ED2DD14697E85AA849";
    attribute INIT_1F of inst : label is "9B7D10AF3162C43B58B079E081E1343F7511881C767101C72AC51C7FCE3E17EE";
    attribute INIT_20 of inst : label is "85CCDACA749B28E228A80069219E386114427139562C722E86191D0C311185B6";
    attribute INIT_21 of inst : label is "C03FFFF07FFFFFCF003FFFC3C03FC1C03FFFF07FFFFFCF003FFFC3C01202A8AA";
    attribute INIT_22 of inst : label is "3C7EFFFFFFFFEFE7C38100000007EDDFFFDE0402FDBE07FC153D3F820E9E9F41";
    attribute INIT_23 of inst : label is "40404B20A282890000000080E0F1FBFFFFFFFF9FFFFFEFE7C381000000001018";
    attribute INIT_24 of inst : label is "B41425118D0028D08216D00A90F31785C44FD9F2E21FB2026DA8041546C78C5B";
    attribute INIT_25 of inst : label is "25AD35A90865C01B100E0108A24B642005AD130008040000276BDB5B0276D6C1";
    attribute INIT_26 of inst : label is "10070D055EA915A05D17225E0122CF8B57235305D234C0560249004DEC15827A";
    attribute INIT_27 of inst : label is "C639C71E1E0FC0000007E0F0F1C738C631CE38E3C3E07FFFFFFC0F878E38E718";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "CA35D03FBAB8ACDF42EC5411F9C7BF8A003D55804AA64304308A28244A00D94A";
    attribute INIT_01 of inst : label is "0EC21B6A3BB43082340D8660AD304695C50035D8134084412000302AB03EEC5E";
    attribute INIT_02 of inst : label is "6DF241475A3769C0866323A2200290A03D113A0427410000003B5AD547D0D2A8";
    attribute INIT_03 of inst : label is "1E674CE264A67C866E83A252810047FE560CAC0111034020F212C20828211984";
    attribute INIT_04 of inst : label is "20E61573BA02111071A38FAD898F8255812F424DC4081B3265459919511A48DD";
    attribute INIT_05 of inst : label is "082CA30BBA7C869991021BC24E004222A61A20B0C2375B126DB46B1067AA5350";
    attribute INIT_06 of inst : label is "CAB95592FF67BF3CB024AAEAFAAF2528336403272708000E32208052D4D24000";
    attribute INIT_07 of inst : label is "1F38DF491E7F1DCF7FE7BFBFF3C0E5714C3400E00E42A0135B0694C284468115";
    attribute INIT_08 of inst : label is "1000040605053F20C9F984A66DB76DB11A084810A101001658DDD5CE531F0420";
    attribute INIT_09 of inst : label is "DBF70F90B5B770F90B49906E491639392E3F5C433A7971641FF0332D0020000C";
    attribute INIT_0A of inst : label is "11A39007E17E88C5054E8400285008069249289F9B7A19FDD64B47DCFF8DF9F9";
    attribute INIT_0B of inst : label is "EFFDC10EF822C9072E091BEA9FB4BFB0081C46456862B74EA022FDA5A6A4CEDC";
    attribute INIT_0C of inst : label is "171300523E777E97830290452C8013403812D16BDDEC67E7FCFCFCB7EE0877DC";
    attribute INIT_0D of inst : label is "C2DB73061FE2C4609E0602231404A10095DC773FFEFD8104B158500E8E4CAB49";
    attribute INIT_0E of inst : label is "884BDE3FE9FB09000074EA487BB7DF917C16542B7BFBFFF9825A8EA010E29D47";
    attribute INIT_0F of inst : label is "007DD4C07FDBE5FBBD8C7CE7FFDF81DA9620FF3FFEFC0ED4B107CBF03BFFF6A5";
    attribute INIT_10 of inst : label is "19009A0B815DEE3188A6D126C936124F2480262AF77B190066037E9F2AF77B19";
    attribute INIT_11 of inst : label is "BEF5FCEEFD6E9B6D7BF7C08D1F0553FDFBE0412C870C28402820001EE8DBFE16";
    attribute INIT_12 of inst : label is "59A01A944CB5FE8A98B1D52D482FEF12A07EEEFA9E4D3497269A4BC12EF6669D";
    attribute INIT_13 of inst : label is "40394571F1020840024481212C2A083A4D96C9E8162253BA463140AC59463583";
    attribute INIT_14 of inst : label is "7F6144ABF482D24824045A07476C9249239C27BCA8F8ADF322B16924BC000514";
    attribute INIT_15 of inst : label is "7E0003FD3C0007FA78000FF4FA07FE70003FF38001FF9C000FFCE0007E014000";
    attribute INIT_16 of inst : label is "4D03A625DB2492492DBE8040DC3280238E0910226A6784495B9FC964DB122AC2";
    attribute INIT_17 of inst : label is "C43400F610D64EA2A1B450834A16008C633E62E1EB37C0758BDE603DC9F6CFD4";
    attribute INIT_18 of inst : label is "511031114A25FAF009108F58AFC8FC0768892FD04ADCFF15150364A8B1765847";
    attribute INIT_19 of inst : label is "55D5551DDD9B6D7F69A5CFD34800D34A87EFB2C813803B1D8E8743A1D8E94111";
    attribute INIT_1A of inst : label is "638389D237208ED07C6342A9012FE42420D4540D9249258B86BD5555D5554F55";
    attribute INIT_1B of inst : label is "0E402AB0F070116A189AC28427200000000000000000000000014D3F83BC18A7";
    attribute INIT_1C of inst : label is "06C3F4EA438B10FCB174138FC2EF399A733D26918118906046046226DB9B6C63";
    attribute INIT_1D of inst : label is "736D8CF9716761500AC3A3AAB88BA82B20A10AA2BF9B3965708AE0A615289A02";
    attribute INIT_1E of inst : label is "012E07A1040400400FEE4E0AAF2C4346B382A031B61404C4691940849CDA8CDB";
    attribute INIT_1F of inst : label is "620311AC31B281251040F06003C1B4676E858A30B7E123FFCCC41E4804724DBA";
    attribute INIT_20 of inst : label is "060F1CECA1BA6AC6A4A91065271A9249D4833399DA9D452A823255046AB08C1B";
    attribute INIT_21 of inst : label is "003FFFCFC03FFFC0C03FFFFFFFFFC0003FFFCFC03FFFC0C03FFFFFFFD082AA80";
    attribute INIT_22 of inst : label is "C381000000000000000000000005491FFFD0055554AAA7FFEBFFFFFDFFFFFF40";
    attribute INIT_23 of inst : label is "6060C10C1020030000000000000000000000005FFFFFFFFFFFFFFFFFFFFFEFEF";
    attribute INIT_24 of inst : label is "CC1A252B5D1479C433B3D0C6D0220FD0C600D9E86301B1146BFE659DEE07CF43";
    attribute INIT_25 of inst : label is "5B8E9B941223848D1B44012224125A8405E5166209A00124A0681BCA2A06F28A";
    attribute INIT_26 of inst : label is "E007EDBD1445066A202A7D4F157A89395923730144AA7CAFE54600B4BC28E526";
    attribute INIT_27 of inst : label is "F83E07E01FF0000000001FF00FC0F83E0FC1F81FC01FFFFFFFFFF007F03F07E0";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "60CA0A0C0AB0D360D2EE069180934040401DDE262FEFAE5604D5D636154E932B";
    attribute INIT_01 of inst : label is "16AF1F7F373E6CD096C8776A85904E4A6AA85B4EA82C800024117916B4A15431";
    attribute INIT_02 of inst : label is "36A372484B2A52820309DEB12003D4203C8069370D2D0000000916B5E7400BFA";
    attribute INIT_03 of inst : label is "18750EAE893A5405CD1230C66C782C507654ECA030525B2C0D91101008034904";
    attribute INIT_04 of inst : label is "C352CB349A0AD9123CA613989A986F487D254CE54FF949A2EF4CD17BD300A2DD";
    attribute INIT_05 of inst : label is "0EB6A90AA34E92D9B3FA49D21A435B2312CA3D965211796C48495312275222A4";
    attribute INIT_06 of inst : label is "1F21E61F92533E2B7615D3D4F53EDC3E1139484D448B136762A3C07291966E73";
    attribute INIT_07 of inst : label is "B0124CFF81E4220FAFE15FC7F0E93659C412002002865FABC8B2B456945D9839";
    attribute INIT_08 of inst : label is "4515059419257F23CBF99C66C9244922561C87D2A77D7294F18F3DC4F430DEA2";
    attribute INIT_09 of inst : label is "8B24E05690624E05691302D9B036A9A98C3658533A4AADE592A002502AAAAB69";
    attribute INIT_0A of inst : label is "11315726C95406EE16AD04AA0C65967292492DE91550116D96424CB9CD1AB398";
    attribute INIT_0B of inst : label is "C4E93D903003891A944951598929492A312C46454132F61C0282494244A75520";
    attribute INIT_0C of inst : label is "B6D764652202C2B4A4E32CAD2928620271129148190D22CE6959CC9649EC8199";
    attribute INIT_0D of inst : label is "E9241BDFED43B56C5D96181BB844A99945DA2225B4807D44A6043FC26F41B489";
    attribute INIT_0E of inst : label is "B81A9C522C92AB000071E07AE16FCD857C97742B3D90F6FDEF5FBDE470C23804";
    attribute INIT_0F of inst : label is "5058FEF65DAF044321A47DE5A6BFDAD7B6E0FF2D35FED6BDB7058F6B51A625ED";
    attribute INIT_10 of inst : label is "7AA8A50D6D557410BC934C9A24D1124B2728392206434A5077B2ED382206434A";
    attribute INIT_11 of inst : label is "173484058D24B64ACE483E9010DDBE67241F4A5254A81240282000294DBC6D7D";
    attribute INIT_12 of inst : label is "E6F642A16A2A444AD2B545A15035F263ED25BB4FA3FBEFA9FDF7D437AA42030E";
    attribute INIT_13 of inst : label is "482D654181443B554A54892932AAE4361B8DC4D87EE0D7F60D3BC5BD6D521482";
    attribute INIT_14 of inst : label is "36080802C1208165B65043498324925931B87B1FB0095227D3F76924A0000D96";
    attribute INIT_15 of inst : label is "263181814C63030298C4060531E17E139C1BF09CE0DF84E606FC263037F84420";
    attribute INIT_16 of inst : label is "01A44024C924964924C5C6F04B77D10940C803222803644B4A8AC924CC132A00";
    attribute INIT_17 of inst : label is "896E6CCB22524FEFE49E24B28A129A92880889185908203440211C407908200D";
    attribute INIT_18 of inst : label is "593805194E256139C9A4A0806919C820C8892B52CA54561FBFA924A899424001";
    attribute INIT_19 of inst : label is "0080003FDDBF6F5F9F7CD73EF940BEFAA67DF0AE94492994CA6512894CA74173";
    attribute INIT_1A of inst : label is "01B220D66A8C4062583172401B40D0033CFEFEA4924B24D033A8000080000A00";
    attribute INIT_1B of inst : label is "9DCCAB76B3721954D3104AA52424000000000000000000000000100CA4E52243";
    attribute INIT_1C of inst : label is "E59961C06A4F134A00A80175AD5C1302266807FD87387163CE3C2256DB5B6CC2";
    attribute INIT_1D of inst : label is "4A49106AADE5D3C84A52A500922122A1AAABA2A0880835E554CD5AE49528B664";
    attribute INIT_1E of inst : label is "03AE52A50404004002028717AB6DC21405B2A500ED0300833FD1428A1E951292";
    attribute INIT_1F of inst : label is "9AC31352A6E28552A7B494E403C3352E78961000A70643FFD16594F7DC742DE0";
    attribute INIT_20 of inst : label is "7C0FE0F0C12C4884AF5B315AF152BAEBA904063332BD8770B29361652AB4A4D7";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000007D55555";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000D554FF000000000000000000000000000";
    attribute INIT_23 of inst : label is "41DC904905241600000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "B9960D2F350089732F5D501295266FAF45C0D3F7A381A41D695299744B8F9AF3";
    attribute INIT_25 of inst : label is "16BD96A61AF186B9592401160926815405B51EE0C9A401B6AD6B5B6B2AD6DACB";
    attribute INIT_26 of inst : label is "A0076082BFAEA4E402C03A5C63657968522A1A9A56A6402001408C2C831A0180";
    attribute INIT_27 of inst : label is "FFC007FFE00000000000000FFFC007FE003FF8003FFFFFFFFFFFFFF8003FF800";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "49A51198103130408C4C6D4C813D000980244FB37AB36EDA5B2BEE626B7B2418";
    attribute INIT_01 of inst : label is "9F827B67F11F625B4A24932432486D33FD5A791F44B64B6DB25C14BE12204490";
    attribute INIT_02 of inst : label is "80625A282FE2C108C4942A0480064398B2456C10AD840000002C9390CD0126AE";
    attribute INIT_03 of inst : label is "94C19833924B160D800A0063D4CFBD5646148C20E1293892104868E385B9A74F";
    attribute INIT_04 of inst : label is "205965DFE80844C1C26A5FAAA8DA07F3C0D9A150A43CA407452E03114B69E6DA";
    attribute INIT_05 of inst : label is "0F8E14F06C6E1922441024195B0108985823CC69292206372CFE6441D3299253";
    attribute INIT_06 of inst : label is "678EF2EF3F6BE518180678BE2F95F3C2E482A92EE68C31CEA143D47C55D792FD";
    attribute INIT_07 of inst : label is "7027B480042409F05005E03803A30D34526DFCBFCA778080379D47A9478440FC";
    attribute INIT_08 of inst : label is "5050508724D3F620DFB18438249724B9B26B3C80F9802D6D5DBD58D551B40F67";
    attribute INIT_09 of inst : label is "E1FE1F82323FE1F82321D96CD8F1F171365B6F088767601009F6DCAA0000010D";
    attribute INIT_0A of inst : label is "1BB982D17C3EF381DDE27401290861AC6D249A7F8A7B8CEC92D017CF7FC75EFB";
    attribute INIT_0B of inst : label is "6BFF808FDCBE861B972D9CCC1FBABFB1C8533131776C3B366EC9FD9FE23047FA";
    attribute INIT_0C of inst : label is "420181081ADDED4C81084310AE547126381ADE2B65B2957BFFAF7DC3FC047EEF";
    attribute INIT_0D of inst : label is "EFFA530673F880701C0623CE077214261C44551E7FDF8812B982590B3827EFE4";
    attribute INIT_0E of inst : label is "C827EB7F7BFB0C0000B3673BEEFD7FD17D471493FBB2F659925ACCB791686CD2";
    attribute INIT_0F of inst : label is "A83BFCC82BE3976CB6522F73FFD7F2F287205B9FFEBF97943902E2FE5FFEFCA1";
    attribute INIT_10 of inst : label is "18DA690F86307E620E5822C11608C92690541CBAD96CA4A826415F5CBAD96CA4";
    attribute INIT_11 of inst : label is "EE4B15BBD2D25B6DDB66C402A4037BADB36206AB26CE4D003FFFFFCDB20D2C1D";
    attribute INIT_12 of inst : label is "048010CA1805016084385108663E2F92B2D20A020900000C80000503C7898C7C";
    attribute INIT_13 of inst : label is "0029040C8C41924069162D0D94E667924924D349920248922573448B1C29E301";
    attribute INIT_14 of inst : label is "5800000F00139C106D0B251938DB69248C07657E636FAD89B49924920C000411";
    attribute INIT_15 of inst : label is "B8000280D0000501A0000A0340058050002C0280016014000B00A00059F94000";
    attribute INIT_16 of inst : label is "B28C9B9236DA4924921C8D78C810A414362404998007132430F1A4DB31C8C125";
    attribute INIT_17 of inst : label is "12248242492DB2B2B2448A0861E868400028000144800053200000014400001C";
    attribute INIT_18 of inst : label is "338889E42190CCC6A41A1000F966CB8A46648669218788759524DB0F661B24BB";
    attribute INIT_19 of inst : label is "0080005999DB6C558003CF0004420000B2492A08C1A08442211088442A150C19";
    attribute INIT_1A of inst : label is "838801F722D2170D31CC4934C43399C08256549B6D24920D88A8000080000A00";
    attribute INIT_1B of inst : label is "6DA002643A351ECB1C96E0D290D0000000000000000000000002002C81A40907";
    attribute INIT_1C of inst : label is "42D1B3672EFE19FE5CBA09F7F96AD98077ED2693211210C844840D224B892E5E";
    attribute INIT_1D of inst : label is "7125CB8760104060A5A85100100900090009080A880970101226C011418F5101";
    attribute INIT_1E of inst : label is "990BAC510404004006901F728F0E4B3649D63DD7372A82F3793084232C5ACC49";
    attribute INIT_1F of inst : label is "2C82192B39A1405DCA8C4E30A98129C57108608E1700800037186660092D39A2";
    attribute INIT_20 of inst : label is "AFF000FF04BD62E2329C437DA09E4924967A4A00164870AE89481D12989A5232";
    attribute INIT_21 of inst : label is "000000000000000000000000000000000000000000000000000000000280002A";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000D554FF000000003FFFEEEEFFFFF777700";
    attribute INIT_23 of inst : label is "004AC92C92B24A00000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "8C1224991412440C3B1142488137D8248400CE1243019C37251021DC210B824B";
    attribute INIT_25 of inst : label is "5C03481128ADCA2C2C9201C896C9252004A41242148004920721C94820725208";
    attribute INIT_26 of inst : label is "0007907815501D70C000788C2932A56B30CB3BC5521D00B0073200E2002C0700";
    attribute INIT_27 of inst : label is "FFFFF8000000000000000000003FFFFE000007FFFFFFFFFFFFFFFFFFFFC00000";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "00A510B83020B00184480080801500C080008FA230015ED66901C74121620011";
    attribute INIT_01 of inst : label is "E9844927911E445B8242000221002832B807A8118DB2496492CA22BE02200010";
    attribute INIT_02 of inst : label is "C96093080360C180421821080006039AA0554001A80000000038918049200405";
    attribute INIT_03 of inst : label is "98C218439254280CA50E02313183A9124210842060313900088000C304B0C34A";
    attribute INIT_04 of inst : label is "20513D5BA9F008004448DE222050031141C88100C000C407C2640330996B2C4A";
    attribute INIT_05 of inst : label is "0D1818502A2950952A011299508001005041A022B5332A13642736A049295252";
    attribute INIT_06 of inst : label is "778EF2EF0932A518200478BE2F95F0A8A0522809C0803549E40314645554A175";
    attribute INIT_07 of inst : label is "30029400002104000003000000E1093460A5003002348018528506B1028C88FC";
    attribute INIT_08 of inst : label is "4054408304E26A01535088184DB26D91F02114084A0005A90528405100A00647";
    attribute INIT_09 of inst : label is "64920481661920481664DB244AA2DBDBB2C924000726204009965EA800200105";
    attribute INIT_0A of inst : label is "EA7080512832E080D0467000190A2884248040048C4B8CB9C64012653CE64A7A";
    attribute INIT_0B of inst : label is "23C480424CB99019522DCCC2049AA49B887A202135342962C4CB24D922208893";
    attribute INIT_0C of inst : label is "8200010A1AB5DD0C00884140A6457166A81A4A2AD56B5129E7253D4924021265";
    attribute INIT_0D of inst : label is "8C901204713180401404038203681832188C1112624480229180300208210250";
    attribute INIT_0E of inst : label is "88666B494249880000962C1BE22564D135035F1990A0A659024A8CB31130C5A2";
    attribute INIT_0F of inst : label is "8A0A7C802B62B35AAD6A25209256D2729220490492B69394910242DA4C929CA4";
    attribute INIT_10 of inst : label is "108C608C823072420C5862C31618809642451D9AB55AD48A24015B159AB55AD4";
    attribute INIT_11 of inst : label is "AEE9156BBA5A4927D1224042800359E8912026AB72662E803FFFFFC0020D0419";
    attribute INIT_12 of inst : label is "6282108214254560C424518842323910035240900992490CC9248401C689857D";
    attribute INIT_13 of inst : label is "0828001888410200401028881484021108140140B40000A00452000A3030A179";
    attribute INIT_14 of inst : label is "180000070000B80001092F08104924801803457807270880A8A0024804000802";
    attribute INIT_15 of inst : label is "9800008050000100A000020140039E10000CF08000678400033C200019F84000";
    attribute INIT_16 of inst : label is "97840B0012492000004C01898822025832440D1B00032280105110491581416C";
    attribute INIT_17 of inst : label is "122004400024900000091810C1603040000800004080001680000000C000000C";
    attribute INIT_18 of inst : label is "121808A801408DE2109C100039634B016050042010828860000049052A092D93";
    attribute INIT_19 of inst : label is "0080004888C924558002850000400000A2492208801004020100804028142820";
    attribute INIT_1A of inst : label is "809000E42080122E215D5170C83799D1040000092490004C90A8000080000A00";
    attribute INIT_1B of inst : label is "3484036423341ACA488280E308C8000000000000000000000002001C00200501";
    attribute INIT_1C of inst : label is "0270962C0E5485250C93E8B3692AD16044C581A3221228C884881416D95B645E";
    attribute INIT_1D of inst : label is "2B6C8BC620414110D4B0490010010001000100001A4050401044402841057221";
    attribute INIT_1E of inst : label is "8088B449040400400692927299044962C88269C512A0FA324A12004374CAAADB";
    attribute INIT_1F of inst : label is "38C08529916400D8C88C5E4030830145510E300C150203FFF708A460010C3922";
    attribute INIT_20 of inst : label is "07FFFF000495226242900120ACCC000096E24211140830C711880E23100C6072";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000030080200";
    attribute INIT_22 of inst : label is "000000000000000000000000000C003000100400000004000000000000000040";
    attribute INIT_23 of inst : label is "004A800800A00300000000000000000000000010000000000000000000000000";
    attribute INIT_24 of inst : label is "8011001A0000400A09100000C105C82438F006121CE00C3205001058010B0A44";
    attribute INIT_25 of inst : label is "14010001608D58246602008A924B6D2800A01440300400000200814000205001";
    attribute INIT_26 of inst : label is "E0070007EAAABC00C00018CC2012AD41304919854014007001600020000C0100";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
