-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "54292AA049326940A502940A502940A502940A502940A5007E532429B205E993";
    attribute INIT_01 of inst : label is "089B026254A2AE108B0803128C0B4C8AA5128944A251283E67CCF99F33E67CED";
    attribute INIT_02 of inst : label is "9679A953D064EC6F8A80FDCADF72815B0B003001139C89625DEF667791EA3010";
    attribute INIT_03 of inst : label is "C72EEC03973CBBE5CF26F933C9BE5DF26F933C9BE4CF267D1A959F33CD4F679A";
    attribute INIT_04 of inst : label is "307C14072EEC72E6C72EEC72E6C4018CE338CE3272E6C72EEC72E6C72EEC72E6";
    attribute INIT_05 of inst : label is "AA1366CA36423F423642564256452B58D6B7B06185CCBF0DFF1E79F3F43E51E1";
    attribute INIT_06 of inst : label is "2A3BC2CB84296C31658B210B2E94B334A7B0C7D0C7D43E915365FE15602BF017";
    attribute INIT_07 of inst : label is "F2A7973CABE54F22FCE2E82955C041251424BB3DE432ECF790CBB1DE472EC779";
    attribute INIT_08 of inst : label is "DC936572F9C8DB91B07236AE46C2F4CFA3EF4FC1E8FA5CADE54FAEF977EA9E5D";
    attribute INIT_09 of inst : label is "44FA760F0260256400108C7A340217B80A08A5A99B295AA559E82458734D34F2";
    attribute INIT_0A of inst : label is "6CB2084FBD3B50095B324D964B7EB7E8136CEBE58A5A012A20408562F449E8DE";
    attribute INIT_0B of inst : label is "95A49F24B258E0C9FE4103596CC9F37D7A13455E4D8B2C8A93EF56DB0226F932";
    attribute INIT_0C of inst : label is "AD5C95574DCEADB7FB97344C0A2EBBCF56D052405B64093280AFB2049B40D256";
    attribute INIT_0D of inst : label is "9D6D215AE39F3AF3D7000A2148C99367E70A009445178D5E9B9E71EBEB6363FF";
    attribute INIT_0E of inst : label is "BBEF555D36FFAFE14842B999BE7E88B3ADD96B875E7B09E2A1354F445BCFC9D7";
    attribute INIT_0F of inst : label is "2C02212D00B4F15EEB9133A51FA4A3F648639D324F7A37A5FFBFBBB733BFB737";
    attribute INIT_10 of inst : label is "797B45AF3797FE8FF71975FC868C499065970C42188462F018C863FE303B9440";
    attribute INIT_11 of inst : label is "29A56B1AD6DB87FFC30286210C42317C80C67031FF1B4BCEED5E79E79E79E79E";
    attribute INIT_12 of inst : label is "CBB39A9ABF748DF3E04F06F913C9947234549E5EC9E249F89D86FB6656DA495B";
    attribute INIT_13 of inst : label is "7500F9B5F48616B1DF3DF3DF3DF3DF2D1566F2FD70AF72EFD73CBBF54F2AFD7F";
    attribute INIT_14 of inst : label is "9FFFFF6031E7072FF2E54972E5409241FD4B72A540B05739F96E9AFD7C05BFD4";
    attribute INIT_15 of inst : label is "B110E2C4779EF339CC05897AD702B49E0AB402C007E7822483FC4143ECC3ECF4";
    attribute INIT_16 of inst : label is "870EC1E74387E0F3A1C3B47BD0E1FA3DE870ED1EF4387F18D1006115E93F3C61";
    attribute INIT_17 of inst : label is "CBFEAF637ABFDEEF7C054BEADBF71A0E66EFFF67FFBB47BD1C3B47BD0E1F83CE";
    attribute INIT_18 of inst : label is "E55B2A31DB651D6386751C97471EDF9589FD6DE49FFEBFAFFAA52FD677A7D67E";
    attribute INIT_19 of inst : label is "A01B1B368C87352ED3BB5D4BB288922C4B9DCB645CEB4288E72BD5EAF1CF1C68";
    attribute INIT_1A of inst : label is "700007400070080740807008074080731D8CB3B7C20A305AA00CDC46B80E751B";
    attribute INIT_1B of inst : label is "28A8F972CE4CA9E0A8888855555552AAAAAB5531D8CB10000740407004074000";
    attribute INIT_1C of inst : label is "EEE44C913040524BA02488AFB051EA5D095D2E8483F88FA1422802104713A920";
    attribute INIT_1D of inst : label is "8805502014045051010810A00B2450069050A1000A08B9EEFDBBEEFEBBEEFFBB";
    attribute INIT_1E of inst : label is "A08E022F78F61084238424F63BDEF0000340000F3D77EAFE54F2A4F1AF029002";
    attribute INIT_1F of inst : label is "A60C60A026029685AF1C3CDB33633B2983AAB58D9A67210AA6009F9BCC4E6B46";
    attribute INIT_20 of inst : label is "100F1E2C58F1E301E04F5EB01EA4DBB0D58C07A92D58C078136EC048098713C1";
    attribute INIT_21 of inst : label is "622883E28881888A2031146032AF7113D05A37C0A385BE1A88EC0B0A46F86A27";
    attribute INIT_22 of inst : label is "06A20880C45182CAB9444F4168DE028E06F02A03F03C091BC0A89EF147C50F00";
    attribute INIT_23 of inst : label is "E13A8AF7ABC422AB5140F79781058E29C1501500595BC50D143C01A8A2068A22";
    attribute INIT_24 of inst : label is "7684F314A0002ABBCB46A08A3F4A5294A5296CF0889148101425F59EB588486B";
    attribute INIT_25 of inst : label is "9E2CF88CD3D751E2A084D102134F5D478A82132994CA653A79CABF5D9E54F2A5";
    attribute INIT_26 of inst : label is "7F1F1F1F12203AC09D109624E884D3D311E2A08CD002334F4C47888233C19F11";
    attribute INIT_27 of inst : label is "2DF55442B404F8888888888888888888811AB800809090808000009292828359";
    attribute INIT_28 of inst : label is "8849951362B8B62BB8AE2D8AEE2BB8AE2DE568D137D583224F560D5B77D509D5";
    attribute INIT_29 of inst : label is "A00845F80D964F89AC00310AA095B10B4800A04B48713440F2BEAA30DA2F2BCA";
    attribute INIT_2A of inst : label is "522D80AE32FF4FFA3FDAA02916E057197F2BFD5FE940148BF01B2C9FD7FEAFF4";
    attribute INIT_2B of inst : label is "2D806397FA7FD1FED50148B703B3CBF937E8FF6A80845B01D9E5FC8FF47FB542";
    attribute INIT_2C of inst : label is "C0AE72FF4FF27FDA802116E057397FA3F91FED50148B6018E5FC8FE47FB54242";
    attribute INIT_2D of inst : label is "34AD635ADFFE8DF6A00855B01D864FE8DF6A80855B01D864FC8FE4FFB50052AD";
    attribute INIT_2E of inst : label is "A2AC0F445FDA2BF3F69C3C9C9C9C9636229D769C369C369C22377C36969C369C";
    attribute INIT_2F of inst : label is "D2BCD95FB1DF2A797281B2EC82F10842485780A092AD2B6BD67B4BEC8B466E67";
    attribute INIT_30 of inst : label is "7A6811111BBBBB11116C7B4B6365B18F6918D91B21ED2C86CB211ED22364579E";
    attribute INIT_31 of inst : label is "3232321210327272321210327272321210327A7A72121032723A7212103A7A7A";
    attribute INIT_32 of inst : label is "0A0D64164825CE4A08904AB2E2658070E6700320A9882C320A92612A95521032";
    attribute INIT_33 of inst : label is "99493300361906B92725001120F927995801912506A98D411A0C02A926233CF0";
    attribute INIT_34 of inst : label is "950080192C913874173CCE4005C03CF0061C93D925F33801D06B92725001120E";
    attribute INIT_35 of inst : label is "E5DF0EFDCE261095D8904A0289082D2C6D093012901412D204A862B120905B2D";
    attribute INIT_36 of inst : label is "B07A67D17E99E5CF2E7953C99E4DF267977CB9E5DF2AF977CBBE5DF2E7977CB9";
    attribute INIT_37 of inst : label is "D5AD55555288894925DA872C0000BFFFF5289575A9D500C5801EA6B1287D33E8";
    attribute INIT_38 of inst : label is "A1942650104FEB12F46D1A368E34D4C00017FFFC895552555155235595D63155";
    attribute INIT_39 of inst : label is "5E9A5FA695FAEFBE7BE38E39E39E3EABC23C6442A74E9D30048480102FA3A38A";
    attribute INIT_3A of inst : label is "4D14D14EE36F244B5C8638DBC913DBFBC913DFE9BFBC913FCC07FBD2B5A528CF";
    attribute INIT_3B of inst : label is "53453453515515515515515515515515515515515514515514514D14514D14D1";
    attribute INIT_3C of inst : label is "6DE4A45152802200000220020254554554554554554514554514534514534534";
    attribute INIT_3D of inst : label is "555555555555555555555555555555555454505055552B58D6B659215D611209";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555553F00";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "83F2E41E8666A5D997665D997665D997665D997665D99764C0634CB1865D9187";
    attribute INIT_01 of inst : label is "64732666DA46F64D9D2B3727FCD86AEEEE7F3B9FCEE7F3284D08A1342284D09C";
    attribute INIT_02 of inst : label is "077D90591A61BC801782769404A6AA333822F2CD9CA19A968779CECE7B467639";
    attribute INIT_03 of inst : label is "DA5C0D992E49704B825C92E49704B925C92E49704B825C96C43804BBEC8477D9";
    attribute INIT_04 of inst : label is "11A32E5A5C8DA5C8DA5C0DA5C0DD97C0701C0700A5C8DA5C0DA5C0DA5C8DA5C8";
    attribute INIT_05 of inst : label is "3E5A3400A008A908A008E008E00E4A40A6DEB2ED8FF89D40E820820C089B74F3";
    attribute INIT_06 of inst : label is "D0A4080096624888484244424B0021ED8B02236223611B22F463FE9A49D2F46A";
    attribute INIT_07 of inst : label is "07403801D00A024E060E019A3C1595E9B50B4DC6898413886F34DE689C413086";
    attribute INIT_08 of inst : label is "8165975602B7016C162DC265B0494B82D805B058B70969525A02D092809400E9";
    attribute INIT_09 of inst : label is "AA25087AEB4DE8D2FB62CCAD40DF5AD25E646D1CD01AD7EBC4BD6AC1CD92D9C5";
    attribute INIT_0A of inst : label is "4424B3D0D2809B5AD005965FD91B1122C9005EEC12136F47968B17644A00B525";
    attribute INIT_0B of inst : label is "CB8D456A76B1CC1B4192CEBB5ADA0E12A174A6C0B641092CF434A82B676B825B";
    attribute INIT_0C of inst : label is "07AC255DF20278E28D280AD0BE5B8034A02976A4F009645BE4F805B26CF226B5";
    attribute INIT_0D of inst : label is "00BDD591C52D64800B72F145B5863C31012E5F628EAD27AC258816CCCC444400";
    attribute INIT_0E of inst : label is "45F19577C83F9FE5E5E4D890A4B5D74CF2E2471C9005166712CDB328E6968324";
    attribute INIT_0F of inst : label is "C9991B582208F27E8723522C448788DAD577FF16D394C34AC0044440048CC88C";
    attribute INIT_10 of inst : label is "0650B3A2D12803404A49FCA925AAE50143343D8A7B91EE387BFD6FFEDCE0066C";
    attribute INIT_11 of inst : label is "1AC94814DBE99296AB8F1EC53DC8F709C3DFA6B7FF6C949E43E1061061061061";
    attribute INIT_12 of inst : label is "94202D075C0125440E005403A01C06AD0A69A5A15A48127919703A118416D610";
    attribute INIT_13 of inst : label is "C3B303CA965E4E7220830C20830C208ACC122501C678ADC13809445A82D09680";
    attribute INIT_14 of inst : label is "0FFFFC147368487FEB0DA5EB0DA65F23FDA5EB4DA65D2252074B0492A0B10429";
    attribute INIT_15 of inst : label is "922A04489BB17421882C0DEBDB66F64C193616025E4A447247FD2589C009C029";
    attribute INIT_16 of inst : label is "15A81E898AD40F44C56A43A062B521D0315A80E818AD403CF224F33C2B820102";
    attribute INIT_17 of inst : label is "5CF45745F35EAEBEB8005BAF7D53E4E94896FFC97FAC7A2656A47A262B523D13";
    attribute INIT_18 of inst : label is "161133303E2602D35818021780BFAFFE14001B50301FDF03FF8A5700FC4BD906";
    attribute INIT_19 of inst : label is "C01EA8BA0A8A4A9A73DEDE16849409208D34CA242AF1200D00B21B0D80248260";
    attribute INIT_1A of inst : label is "7400070000700C074080740C0700807618CE18F3800400E9400A9A0034836C03";
    attribute INIT_1B of inst : label is "F9F62C0590B96F0075F5F50CCCCCCCCCCCCC66418CE1A4040700407000074040";
    attribute INIT_1C of inst : label is "800EC183108C8F069EDFC55AB32B87B99B801A7B56022A5FA7EF71A3E9E028FA";
    attribute INIT_1D of inst : label is "CE9F73F3DA6C7BA21E17C93ABEFEE246ABFBEBEBFE3DF4801A00801902801902";
    attribute INIT_1E of inst : label is "77D1D03AC3EE318C6696E8EE7EB586DB6FDB6DB856E0B720B905CA0F1AEDEF15";
    attribute INIT_1F of inst : label is "FDFDEAEAD8545B9DFFB9F328B892130101F01C945C2C05BFEA49C0F18481C0E2";
    attribute INIT_20 of inst : label is "FFD1B37EFD9A3D6B5C91A3D6B5493BB3EBD4AD7A5FBF4AD5A4EECD2DAF7A6D37";
    attribute INIT_21 of inst : label is "A5C55C95457AB72DCF56E28F445C5AB4BFA1483C5DFE41E577D7F5FD2907B5EE";
    attribute INIT_22 of inst : label is "EADC973D5B9A3F1175EB92BE8D21717BF90BF5EF7FDFD5A42F57B9C4BB2BD2BE";
    attribute INIT_23 of inst : label is "125595D55AB1A95A14BDD5754F5ABC55E92B5F36F22712FEAA4BFAB7355F5735";
    attribute INIT_24 of inst : label is "CFCE0D6784926F3FE0E277D0A8BDF18C6318D5A93D3B3EA54B4FB0655159D3C6";
    attribute INIT_25 of inst : label is "7373C57384A9E25C557BBAD5EE12A7897355EE4422110886029704B140B905CB";
    attribute INIT_26 of inst : label is "EF5F5F5F51335DEFFBAFFF5FDD7F94BFEA54557FBBD5FE52FFA95155FE6A78AE";
    attribute INIT_27 of inst : label is "B6DF8A9BD9A9D0000000000000000000088372005040405050000050504040F3";
    attribute INIT_28 of inst : label is "329248A40701C07009C0701C027009C075DFAD52577E35C4ACFA546CEE189218";
    attribute INIT_29 of inst : label is "56BDA107E271B03370001B35737F067E249BEDB4ACD20AB167D9F1456D36FD9F";
    attribute INIT_2A of inst : label is "ED0A3F51CD85A02D4A457AFE851FA8E6C25C16E522ADFB421FC4E3612C0B7291";
    attribute INIT_2B of inst : label is "0A3F9A6C25012A522BDFF429F54E3616A0952915EFFA14FAA71B0B405A948AF5";
    attribute INIT_2C of inst : label is "7D110D84A82D0A457AFE851E8886C2D412A522BD7B428FE69B09504A948AF7ED";
    attribute INIT_2D of inst : label is "3929029B780B409156BDA14FA271B0B409156BDA14FA271B09405A148AF5FD0A";
    attribute INIT_2E of inst : label is "F35E3FE6B44380809DC89DC89DC89D629DC897C837623D6297C83DC897C837C8";
    attribute INIT_2F of inst : label is "A2EEA97662805882C5CC5819378BBD6579A52C7FEFFB9CD68080001AD6C9157F";
    attribute INIT_30 of inst : label is "F2DEBEBEA1414014147AA28BDAA5EA145122A922A28A2A954AA2A8A25AA4BDA8";
    attribute INIT_31 of inst : label is "F2F2F2C24032B2BABA824032B2BABA824032B2F2FA824032B2F2FA824032F2F2";
    attribute INIT_32 of inst : label is "D100EB2F2482E3267A4905EF9904369C620CF012278493012279E0B319824032";
    attribute INIT_33 of inst : label is "7F2CB5EF9984905CF1933CF49235D78833EF426994CE2DEFDB29A45CB18112D6";
    attribute INIT_34 of inst : label is "DB6D24BFF6DF061246BC439F78DA5AF2C185352EFAD106784905CF1933CF4923";
    attribute INIT_35 of inst : label is "4B807C1297E969DABDBF2F2D3EBF9B9AFA5F5F59FB2BED3D6FD2BDDF6D24FFF6";
    attribute INIT_36 of inst : label is "0BAD41684B420B805C82C09424A025012C49624B005882E01724B825C12E4972";
    attribute INIT_37 of inst : label is "7FFFFFFBF7FBBBBBFDD64AAC0000BFFFF1FEFE7060BA678C71E1926BFFD684B4";
    attribute INIT_38 of inst : label is "672E1EB079A0943D4152C0A9628452C00017FFFDBBF9FFDFFFFFF7FFBBFFBFFF";
    attribute INIT_39 of inst : label is "76104D269B6DA69A6DA61A61861A4350154259BD143850EBFB7FEF6F5058581D";
    attribute INIT_3A of inst : label is "EBAE3AE270EC7E2370E30E3B1F89FB3F0F8992D9B3F0F80B99C19080200802A6";
    attribute INIT_3B of inst : label is "BAEB8EB81AEBAE3AEBAE3AEBAE3AE3AEBAEBAEBAEBAE3AEBAE3AEBAE3AEBAE3A";
    attribute INIT_3C of inst : label is "5DB686593602020000020200000EB8EB8EBAEB8EBAEB8EBAEB8EBAEB8EBAEB8E";
    attribute INIT_3D of inst : label is "555555555555555555555555555555555555555555564A40A6DFD5018E39E3CE";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555557F29";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "55E6CAAE3745B376CDDB376CDDB376CDDB376CDDB376CDD87C690CE4A6749C86";
    attribute INIT_01 of inst : label is "932A05409324A8614A9B8215085692F137D3E9F6FB7D3E5FA3F47EAFD5FA3F51";
    attribute INIT_02 of inst : label is "C451384F0321C8628501B7F50EF4381A1699A7BB752D56B58A50A8B5A2FA68D3";
    attribute INIT_03 of inst : label is "B7D0AB33EA1F40FA87D0BEA5F42EA87D4BE85F52FA17503A84A80EA289E24513";
    attribute INIT_04 of inst : label is "00150A77D0AB7D0AB7D0AB7D0AB11C1C0701C070FD02B7D02B7D02B7D0AB7D0A";
    attribute INIT_05 of inst : label is "462475B2A002A902A002A902E0021182854620AD26FA0AE1A30EBF76ED9A7051";
    attribute INIT_06 of inst : label is "92AD821218AA482A9154815004454892A020AA40EA454010AD4D54A5CA6EADB5";
    attribute INIT_07 of inst : label is "7DD3EE9F74FBB745AE45B8F61B060658210C922DA45B6C24906DB29361248B6D";
    attribute INIT_08 of inst : label is "DE924D25ABF42BEA527D4A4FA14EEA97D02FA049F4099F50FA07D03EA1F42FBA";
    attribute INIT_09 of inst : label is "A07508D74C3A5B5D199328754260677A153BAB0DD6D6B55AB7D45AB0F369A4B3";
    attribute INIT_0A of inst : label is "2C24EEB57EA1C216B17A49352B4934932352548B00CED2DAE9DC9842EA85D50E";
    attribute INIT_0B of inst : label is "068B735BD5B8B806BAD30522DC56AD3AA02DE087491B003BAD5FA072D4581D26";
    attribute INIT_0C of inst : label is "A2DB3007DB45010557E81CB4E51D635EA079D5A602F447264F817A23922785AD";
    attribute INIT_0D of inst : label is "E9FA463E7BD2B25D5E832EF8EC070E74593263DDF3BAB2DB3BC22C6666EEEEAA";
    attribute INIT_0E of inst : label is "2B5A001F6D756D5A7A7838400F49DD4E5DB3F9E64BAE3D99E7B0ECDF39E90592";
    attribute INIT_0F of inst : label is "0774C2D49837A680704AC4955242AA48B075CE84B2DA83AAEAAEEAEEEE266662";
    attribute INIT_10 of inst : label is "98833D0A03EA5DD4EF48489D8488CDCB62AC6B4AD6135880D6F05B54E9063DD3";
    attribute INIT_11 of inst : label is "96423050A8E212566889B5856B09AC5516B7D42DAA757352ABA69861A69861A6";
    attribute INIT_12 of inst : label is "F402AD4DB0442C16FB27DD3EEDF740F500096EA816EBB3810560C68051A4B146";
    attribute INIT_13 of inst : label is "28CCEB0D133535A8D34C30C30D34D350F5087D42692CF50BA85D40FA07D4BEA5";
    attribute INIT_14 of inst : label is "064926542815C7554CAE72ACAE732982AA72ACAE7329856A56C443AB44C46F36";
    attribute INIT_15 of inst : label is "398B84E607A8F6A52C0B1B6EB3D3AD0C4CAC058936EF44BCA6A9C60352034001";
    attribute INIT_16 of inst : label is "936747AB49B323D5A4D9D5E8D26CCAF46936657A349B3A907084702B03C015C2";
    attribute INIT_17 of inst : label is "9ECEF6EE99D9EDD3B1150AFE4AF2B6A52DFBAA7DD5365E8D4D995E8D26CE8F56";
    attribute INIT_18 of inst : label is "274EBA7249D724A95686A4314919EC6A1B636C6423D9586C654B6636826F1CDB";
    attribute INIT_19 of inst : label is "A3D8B6140B0174E560B885355F87F18E7E9219DCEC282A6D693ADD6E3244A4E9";
    attribute INIT_1A of inst : label is "780C0780807C08078080780C0780C07B32C75CE8C0021073800B0A0814102820";
    attribute INIT_1B of inst : label is "E9587555BFF352C00A00AA83C3C3C0F0F0F078132C758C0C07C0807C0C078080";
    attribute INIT_1C of inst : label is "F329A54A81C9DC569B6986F6287DE69DCBE55B69B53EA8E98724CAC2A989055C";
    attribute INIT_1D of inst : label is "8A0D51A7B3B6DED76D670E3DD3998384032BAD9993733EF33E4BF33F49F33E49";
    attribute INIT_1E of inst : label is "64EEC116A4F494A53304D8B5252D49249324924FFAE1F62FFB7FCBF6D6CCE6D1";
    attribute INIT_1F of inst : label is "4312931317BF8D9E1AB76EB61CFAD9DD4AE75A5B0AD581335876C7ED462681C0";
    attribute INIT_20 of inst : label is "085AD5AB56A7472DF2DA7472DF2DAAA89D3DB7E368D1DB7C36AAA421C26772B8";
    attribute INIT_21 of inst : label is "EF2D9947ADA3BC87246386E4EF3BB3C7F27365AC71272D69C1A91A466CB5A72D";
    attribute INIT_22 of inst : label is "8EF23C918E0B91BCEECF5F89C59631C09CB1A716A46938B2C61CB5A1E68E1F88";
    attribute INIT_23 of inst : label is "339E17B1C8D0A1C870F1B1B1DB0B5A596A5AD238A796879A3D7E239C96651C96";
    attribute INIT_24 of inst : label is "653676D7DB6DBB8001C064E2A3D3A94A5294B54991A77336F7AB4A7FBB1999A5";
    attribute INIT_25 of inst : label is "2595A9C157E27BF0F9C52CE7155F89EFC1E714F2793C9E453FD70FB17FFB7FCA";
    attribute INIT_26 of inst : label is "D000000003917EB6B53825B5A9C147F273F0F9C52CE7151FC9CFC3E714B6B538";
    attribute INIT_27 of inst : label is "9BEFD6D06D6DB55AA55AA5555AA55AA55331EA000202420242000052124202A2";
    attribute INIT_28 of inst : label is "94FF0DB625C9625C91725897245C91725CFFC5C7F3FF170FCFFCDD36DD0DBF0D";
    attribute INIT_29 of inst : label is "473381E677AB5466EC1048313326CCD5DB6D39DAB098999377FDFB61B7177FFF";
    attribute INIT_2A of inst : label is "8C0F33BD1AAFA8750AD53DCE07B9DE8D57583AE56A8E6703DCEF56ABAC1D72B5";
    attribute INIT_2B of inst : label is "0F73EED57543A856A9EE303DC6F46ABA81D42B54F7181E637A355F50EA15AA7B";
    attribute INIT_2C of inst : label is "31BD9AAEA0750AD53CCE07B8DECD57D03EA56A9E6703DCFBB55D40FA95AA7B9C";
    attribute INIT_2D of inst : label is "88460A15181D50B54F3181EE37A355D50B54F3181EE37A355D50EA15AA799C0F";
    attribute INIT_2E of inst : label is "587032B0ED1BABA1E88882222288228822882822888882222822828828228822";
    attribute INIT_2F of inst : label is "B62CB316A847FDBFE520AAB97B6D99D150D5D84924DAD4B510C8446B679EED89";
    attribute INIT_30 of inst : label is "3C1B154001540015406212DB12CD89425B14B317704B6DC59B7584B6B2CD6584";
    attribute INIT_31 of inst : label is "3C3C3C0C80347474744C80347474744C80347C3C344C80347C3C344C803C3C3C";
    attribute INIT_32 of inst : label is "0160534C011038039C0220554028001D420F3C847AE923C847AAB8BCDE4C803C";
    attribute INIT_33 of inst : label is "89C718D341E020071C01CF380428E2081CD38900020700530004900554111540";
    attribute INIT_34 of inst : label is "96000069249707808D1041E79E09144499E081C71C61079E020071C01CF38042";
    attribute INIT_35 of inst : label is "FB07FDBBD2C2D0564343414325A58081A034161052196B08C2B1AC0200002924";
    attribute INIT_36 of inst : label is "2DF54BAA1D40FB87DCBEC5F50FA07D43EC5F72FB17D83EE1F72FB17DCBEC1F70";
    attribute INIT_37 of inst : label is "AA56AAAEAD6666E6D38485C000003FFFF5E6B70080B2724B69DDB2E8EF7A85D5";
    attribute INIT_38 of inst : label is "92326AC9A99AB89E455342A9A00188000007FFFD76AEADAAAAAADCAA2A298EAA";
    attribute INIT_39 of inst : label is "24DB6994524934D14914D14D34D11F955BBF39CE3A64C9DD1D39A6739068684D";
    attribute INIT_3A of inst : label is "C9DC9DCBC17D5C171462E25F5705CF7747076908F77470F344A26635AD635819";
    attribute INIT_3B of inst : label is "727727727DC9DC9DC1DC9DC9DC1DC1DC9DC1DC9DC1DC9DC1DC9DC9DC9DC9DC9D";
    attribute INIT_3C of inst : label is "244182082180220000022002023F727727707727707727707727727727727727";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555550505555505211828547148211508049";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555552C28";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "D56406AA216F1EAD5EFDEAD5EFDEAD5EFDEAD5EFDEAD5EFC57581ADD2D6C8C0A";
    attribute INIT_01 of inst : label is "FBDF2AE7C3BE2A7DEAD5EF33BC8C98F175FADD7CB65F2D5FEBED7F8FB1FE3ED0";
    attribute INIT_02 of inst : label is "8EEAC8E3030284FA8621F4C7039610113C9BB7BF7B5BBC6B0948CD6371383CE9";
    attribute INIT_03 of inst : label is "FB1C37F58C4C6263931C18C0C6073831C98E4C6263139C9CC08802F75662EEAC";
    attribute INIT_04 of inst : label is "184D0E7B1CBFB1CB7B1CBFB1CB715F8C2318C230B1CBFB1CB7B1CBFB1C37B1C3";
    attribute INIT_05 of inst : label is "606665B22002290220022902200304315555DE47DD5CB84120138A142B74E581";
    attribute INIT_06 of inst : label is "B22902949EA85822011001100C654810A840C80088044070F839FE63865CFBAE";
    attribute INIT_07 of inst : label is "19C8CE06723381771A77182C1667F7F03006D36DB49269B69A6D349349B4DB69";
    attribute INIT_08 of inst : label is "FC924DE71EC72D8C52B1CA56394D739398B7314AE629EE6063031C98C4C60339";
    attribute INIT_09 of inst : label is "3831CA71EF32B30F85EBCCB9C27D794A1A7BE60D96CC66F3611E72E0726934DF";
    attribute INIT_0A of inst : label is "2900CDE35CC0C3ACE7F249340A002003221B73060C4C95987C2F5E257382E706";
    attribute INIT_0B of inst : label is "FD6E1F30FF18F86FD6A343379F3C6B18E198D0B6594A403378D73033BF337967";
    attribute INIT_0C of inst : label is "FCB73FF30BC76797358E0E60DD04C6D73039B726EFE4CF66CFF7F267B267B739";
    attribute INIT_0D of inst : label is "E867D7CF3C92927D45EBEE78FEC3C760383C79DCF3EFFCB7334E3F27272727BB";
    attribute INIT_0E of inst : label is "F6BAFFCC2EFFF7FF1F1DB0F8724B5D5693633CF24FA79FD9E3F0FECF3C49C493";
    attribute INIT_0F of inst : label is "666CD78C9A2F52B0D56F9E450018A001E29461CF66F242A29FFBBFFBFBBBFBFB";
    attribute INIT_10 of inst : label is "8A892D8E59CE06423952A0C54D980C8B23F8C6EF8DDE34B58D5AB5FE4B5699B3";
    attribute INIT_11 of inst : label is "DC60862AAABBDCECD3BCE376C6AF1B45AC6A95DAFF26D2502B928A28820820A2";
    attribute INIT_12 of inst : label is "C709A9816E8408043281900C846C00B9C10FC7305C2F3005FD30BC9251366144";
    attribute INIT_13 of inst : label is "E4EF1A0B9FC3CAFE5145145144104110B54339C32DA4B9C98E4E6263931818E0";
    attribute INIT_14 of inst : label is "88924C2A1E1901D02E6BBA8E6BAFAFEB07BA8E6BAFADF94AB58C630AE2F4462F";
    attribute INIT_15 of inst : label is "BA99A6EA5694D129490E7F546ED31B3AD5DA873B3529D6AEB7FCF7C240424078";
    attribute INIT_16 of inst : label is "A68F53225347299129A390C894D1E8644A68E432253473CBC3C0A3FE614B0CD3";
    attribute INIT_17 of inst : label is "D642323288C8645193ABE515AC61972E7659FF2CFF974CA99A394CA94D1CA644";
    attribute INIT_18 of inst : label is "4604321288862981C0A128110A086512892DA635014A4AB4293DF25A54BD064C";
    attribute INIT_19 of inst : label is "800AA4100E205180E08A8404548D01000C394884382265684A3090482281A821";
    attribute INIT_1A of inst : label is "3004030040300403004030000300003331C6BA6400000060200E0E0A1C143828";
    attribute INIT_1B of inst : label is "79DC3D05023939C00AAA00003FC03F00FF0180131C6B80040300403004030040";
    attribute INIT_1C of inst : label is "73AD62ED8AFFAF4452CB846CDABB76A570F5104B130E887DC5C6FAAB24B0451A";
    attribute INIT_1D of inst : label is "2B8B632367378CFBCEC76D9DFB9DEB4D1589EA9DB3336C7BB66F73B76F7BB76F";
    attribute INIT_1E of inst : label is "6553C07CE6B2E5395F04F07767B9CD34D3B4D3495CE0E7233119C89DDCCFFCBB";
    attribute INIT_1F of inst : label is "6DA853D3D5A7850AD7CC5DE419D0F1E0A4C13A120806213BF06CA1DDC0C155E0";
    attribute INIT_20 of inst : label is "6B58D1AB568306BD3C48306BD3C4D57A8D1AF4D128D1AF4F135D6AA5E36B74BA";
    attribute INIT_21 of inst : label is "C7D5BC37F5B79FC7F6E3EAD67F369BE26B3D7E977C33F4ADF7619867AFD297E3";
    attribute INIT_22 of inst : label is "DE7F1FDB8FAB59FCDA6F89ECF5FA5DF0CFD297CDA6699EBF4A5F8F78FA6F89ED";
    attribute INIT_23 of inst : label is "03CD5778DC4EBCDC5E6978B8A9E3075D8A2B4BBCDF9DE3E9BE27B71F56F4DFD6";
    attribute INIT_24 of inst : label is "5B7714DF134D39D0F5E0655220F978E6398E66E1B160762C075CF51368F589B3";
    attribute INIT_25 of inst : label is "319263F1E278313C6FF1DCBFC789E0C4F1BFC7F3793CDE4F0AE70639133119CA";
    attribute INIT_26 of inst : label is "B05050707D5566B2ED7EB5966BF5E26A313C6FF5DCBFD789A8C4F1BFD6326C7E";
    attribute INIT_27 of inst : label is "8B34FAFF6FAE7EEBB1144EEEEBB1144EE338D800908080C0C0000090D0C08163";
    attribute INIT_28 of inst : label is "9ACBFA97B5ED7B5ED5735ED7B55CD57B5A34D5BB689356D6F34F5AB7BB9A8B9A";
    attribute INIT_29 of inst : label is "467181E667E2466FF012393FB3F5CDE49E7DB1D7B6C30DE99E65997596996659";
    attribute INIT_2A of inst : label is "9C0F737F52B728390AF139C60799BFA95B181CC5788CE303CCCFC48D8C0E62BC";
    attribute INIT_2B of inst : label is "0F33FA95B101CA5789CE703DC4FC4AD880E52BC4E7381E627E256E507215E273";
    attribute INIT_2C of inst : label is "713F12B628390AF138CE07989F895B901C85789C6703DCFEA56C407215E2739C";
    attribute INIT_2D of inst : label is "8C10C55553EE50BC4E3181E627EA46E50BC4E3181EE27EA46C507215E2719C0F";
    attribute INIT_2E of inst : label is "98613130CC57AB80422228228222282282222222282282882822822222882822";
    attribute INIT_2F of inst : label is "02B0015830191888C5887A111AE9D14150B0B849B6F39CF7906D44CA65FCDD88";
    attribute INIT_30 of inst : label is "2A3A400014000140002A00095004A88001080108300020C00830800210043600";
    attribute INIT_31 of inst : label is "2C2E2C0A10222624200E10222624200E10222A28200E10202A2C260A10282A28";
    attribute INIT_32 of inst : label is "D368D34D0582EB079E0B04D7486D368D020F3C16298483C1629E603F1F8E102E";
    attribute INIT_33 of inst : label is "B95D70F3C1E0B04D74834F34162BAE0834F34160B05D60F3C160B04F3C811DE6";
    attribute INIT_34 of inst : label is "1612096804070792C77C41A69A0B15C249E0B14D34C1079E0B04D74834F34162";
    attribute INIT_35 of inst : label is "6281908A5AC0C0D70B0B0B0BA5A5818184309602D05D6B18C6B1AE9690486020";
    attribute INIT_36 of inst : label is "25B1898C4C623211900CA0E6073839C1C84E427291948C846406283141880C50";
    attribute INIT_37 of inst : label is "2A52AAAAA54222E2D105408000007FFFFE65369AC010BB6E4DA579CCCE58C4C6";
    attribute INIT_38 of inst : label is "1AE5F197CDDB97DCD4534A29A4982000000FFFFE66ECAD2AAEEA942A6629CEAA";
    attribute INIT_39 of inst : label is "749B65B49B6920CA28269A6C36C225F39BCB1AC7B76EDDF91919A6F3BFE9E9EF";
    attribute INIT_3A of inst : label is "40840841BCA8041920026D2A010768300106FBF08300106E0223D8800000041F";
    attribute INIT_3B of inst : label is "1021021088488408488408488408488488488488488488488488408488408408";
    attribute INIT_3C of inst : label is "3041A00040000000000000000062102102122102122122122122102122102102";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555551545555515304315554005010404108";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555550CA1";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "80583C034014AD5AB122448956AD5AB122448956AD5AB122966D1896AC4C76C1";
    attribute INIT_01 of inst : label is "6EC0BC57AAED485932716AB402C258E892090492492090A4548A93526A454897";
    attribute INIT_02 of inst : label is "0410101CEBB0228AD7EBB5873CC724AAB232C6EDDE60129082400188408C266F";
    attribute INIT_03 of inst : label is "9E18C99B4E7A63D31E9CF4C7A73D31E9C74C3A71D30E9870C3288CA080830001";
    attribute INIT_04 of inst : label is "9D59AC5E1849E1849E1841E1841D172A4A02A0A0E18C9E18C9E18C1E18C1E18C";
    attribute INIT_05 of inst : label is "3156B044AB2C86AC8B2CA22CA22858FA38888374099AE942ACA49224591A774A";
    attribute INIT_06 of inst : label is "B4A22C0E165032DA2251165119A93CC948EB288B2889446AE4535546D4F6A2FA";
    attribute INIT_07 of inst : label is "E98F4C7A61D30C50B390B5C2A125A58AB9804160808801104320840928105020";
    attribute INIT_08 of inst : label is "312496D0B387370E62E18C7C3189D31E18DC398B86317873D31E9874E3A61D31";
    attribute INIT_09 of inst : label is "39E985440B448996D572E2E1CD5A5E63542EC95EC102950816020815C496D948";
    attribute INIT_0A of inst : label is "5434991670E72B8214849259950D5042DD0414095411244CB6AB9755D39F873C";
    attribute INIT_0B of inst : label is "3A496C4B10B540194CB268084002C834C6053AF892450426459C31C26009424B";
    attribute INIT_0C of inst : label is "02E13AA60BC49459674C701090D52D9C31C12085AD89CE4B46D6C4E724A32085";
    attribute INIT_0D of inst : label is "8840A49B6DB7B6D14432536ED74376B181264DA6DB1152E03186247666667614";
    attribute INIT_0E of inst : label is "0C08AA982D353D4C8C8D5928E6DC0AA75E036DB6DA269A0DBB40D06DB4DB45B6";
    attribute INIT_0F of inst : label is "C8CBB84077DB0B01AD88584A411B486A16C52900105CEBC8E444404004000440";
    attribute INIT_10 of inst : label is "7146B2E2330E38F1CC4BA131CB772E0B82A5B9CD7399CEEC731E4D556AC8032E";
    attribute INIT_11 of inst : label is "020B1F47112B1B171E1C5CE6B9CCE6796398E726AAB59D93C20CF3CF3CF3CF1C";
    attribute INIT_12 of inst : label is "A61E3000C4D83457D31EB8F4C3A61AE1C7AD2C30C28CC001A22B034120C01483";
    attribute INIT_13 of inst : label is "ECBB63EED6E0E5079E79E79E79E79E6ACA0E61CD06D2E9870E3871D38E9870E3";
    attribute INIT_14 of inst : label is "0649228D473EAC654A8D2F2A8D36F36AA92F2ACD36F17E736459ACB7A0B82CB9";
    attribute INIT_15 of inst : label is "0326660C8BA3764713A12D8B1B64C66F9107D092588E744646AA65AD442D4404";
    attribute INIT_16 of inst : label is "53846BDB29C2B5ED94E15AF6CA70AD7B653846BDB29C22610A7A8BA932010333";
    attribute INIT_17 of inst : label is "B686346298D0E8D3A2BEBEEF34D4938538DBAA6DD536AF6C4E11AF6CA708D7B6";
    attribute INIT_18 of inst : label is "50708164B6104A580928CAAC92B0E8AA1B636F793951516C45493C36AB260CD9";
    attribute INIT_19 of inst : label is "4004108AD1A222591244521081326830730E121A9691080012800A0584A04ACE";
    attribute INIT_1A of inst : label is "0408004080040800408004080040800402004019FBFFFF196011C05280A7054A";
    attribute INIT_1B of inst : label is "094B6E02AD2898400AAAAA00003FFFFF00000040200404080040800408004080";
    attribute INIT_1C of inst : label is "022783265D999B834DB601602733104F30C60D36D0A72B223C519D73B13076D7";
    attribute INIT_1D of inst : label is "64B226424A492927929489D325933249F5AC06796C2EE00A30080A310802310A";
    attribute INIT_1E of inst : label is "333980001125295AC6328AA0F080225B25896C94F4C7861D30E9874C00DEC9A6";
    attribute INIT_1F of inst : label is "9E72925248D6E7CA9AA40A90840A2801481644C8443A0CAC4A496440ACC88E60";
    attribute INIT_20 of inst : label is "085A64C9932B56366CCAB56366CCA206AD58D9B32AD58D9B32881E296A9E4F27";
    attribute INIT_21 of inst : label is "C645E52645CB9946797332F960B28326DCB16814654B40A1952258962D02A641";
    attribute INIT_22 of inst : label is "2E6519E5CCCBE582C84C9B72C5A0D1912D06A640896258B41A192438CA0C9B72";
    attribute INIT_23 of inst : label is "925B1731B8CAE4B8D25D31B1AB230259480A522EA050E321326DCB1917941917";
    attribute INIT_24 of inst : label is "9049442705B245450E60333CAC4F85084A5012292F58ADEB0AEA4A37CA199990";
    attribute INIT_25 of inst : label is "A4D4299526DAB36E699126A6449B6ACDB9A6440904820100A7A63D38ED30E984";
    attribute INIT_26 of inst : label is "14A484A48999669A8532A4D5299526DAB36E699126A6449B6ACDB9A6449AA532";
    attribute INIT_27 of inst : label is "CB76D2D16DAD3FF4411FF00FF4411FF003318A00501000302000004050702002";
    attribute INIT_28 of inst : label is "96DB089605A9605A816A5816A05A81625A76E5AB69DB9696F76C5AB6113ACB3A";
    attribute INIT_29 of inst : label is "3DAD4A24B971750904810064764811152492453C28930329316C5965B69316C5";
    attribute INIT_2A of inst : label is "6A11658BCBAC31E18508D6B528B2C5E5D694F0A2867B5A844972E2EB48785143";
    attribute INIT_2B of inst : label is "51255C5D698F0C2866B5A8449F2F2EB4E78614335AD4A2CF97975873C30A11AD";
    attribute INIT_2C of inst : label is "678BCBAD31E1850CD7B528B3C5E5D61CF0E2846BDA844957175A63C38A11AD6A";
    attribute INIT_2D of inst : label is "8163E8E22018634235EF4224F171758634235EF4A2CF17175A73C30A19AF6A11";
    attribute INIT_2E of inst : label is "1F67F23EC48D80E3888888888888888888888888888888888888888888888888";
    attribute INIT_2F of inst : label is "A442AA21C0869474A2CEDC0C4C22252D33ED20364B421094A4B491303F9BB4B9";
    attribute INIT_30 of inst : label is "2E0180000000000000102A908AA847055272AA70C8AA433550CB0AA46AA8C80A";
    attribute INIT_31 of inst : label is "2E2E2C0800242424240C00242424240800202A2A200C00262E2E2608002E2C2C";
    attribute INIT_32 of inst : label is "080441842110202208422041010080462644108462A11188460829C0600C002C";
    attribute INIT_33 of inst : label is "2B04144108C42204101104108460829910410844220404410844220410133050";
    attribute INIT_34 of inst : label is "4AD96CA592CB23108C14C8820842315088C42304105322084220410110410846";
    attribute INIT_35 of inst : label is "D38E987311594B4A6565656536B69292B2D64AD94B29AD295A5694DACB65AC96";
    attribute INIT_36 of inst : label is "36E98F4E7A63D39E9CF4E7A63D31E98F4E3A71D38E9C74E3A71D38E9874C3A61";
    attribute INIT_37 of inst : label is "FFFFFFFFFFFFFFFFFF105A6000003FFFF775BFA740B833611B3186129CB4C7A7";
    attribute INIT_38 of inst : label is "8E50934A41CB086A894504A280BD1A000007FFFDFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "349B4926D24936DB4DA49249B69218E40EE3A863850A14627272CB5AD020203C";
    attribute INIT_3A of inst : label is "0080880818200001010014080000682010000480820100000009000000084004";
    attribute INIT_3B of inst : label is "0020220208008008008008008008088008008008008008008008008008008088";
    attribute INIT_3C of inst : label is "450E800000212102022303002202002002002002002002002002002002002022";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555505555515058FA3889A01008271A60";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555550C25";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "BC5325E299DC64C993264C9976EDDBB76EDDBB3264C99324F84B28B5945C6D93";
    attribute INIT_01 of inst : label is "264E20C40A70694A1A352A3828A135E6582C161B0D86C3542A8552AA554AA954";
    attribute INIT_02 of inst : label is "10820150CB6488A597B3FC048086A33E31766E64CA1331084802108866462225";
    attribute INIT_03 of inst : label is "181291980B405A02501680B404A02401680B404A02501600B5A810A4900B4920";
    attribute INIT_04 of inst : label is "11012D581291812918129181291D562A8AA288A2012998129981299812998129";
    attribute INIT_05 of inst : label is "944DF00E804E84CE84CEA04EA048807C010083DC1B33E447A324D3AF4D9AFF23";
    attribute INIT_06 of inst : label is "7EA04E0352780CE84F402750213D2EDBE013A133A01D40C2E2D755DABDD5A669";
    attribute INIT_07 of inst : label is "21E10F087843C0544294610138A4A4C4B53124D6D9A597D966965F259ADB7C92";
    attribute INIT_08 of inst : label is "B124978C4204A0094B012960252B02C01600242C0485205802D01280B005843C";
    attribute INIT_09 of inst : label is "24012352490DC4C24D2A78816948484240AED09FC02108068840858905965B88";
    attribute INIT_0A of inst : label is "1C02BB8840B00A310CC4925DBF09F09ADF09D49890836E26126953C4024005A0";
    attribute INIT_0B of inst : label is "5090888408410CBA809A4844297108C090A222D0925700AEE21024063CC4424B";
    attribute INIT_0C of inst : label is "0D29AAA4820A4410040B418EB4C514102C057C758909564B56C484AB24AB3C42";
    attribute INIT_0D of inst : label is "9808849145B6B6D3423A5144809A84F044A549228A140D28AB88524444444440";
    attribute INIT_0E of inst : label is "954CAA9208951544A4A6BAD386D8A014A28A4516DA65104512088228A0DB9DB6";
    attribute INIT_0F of inst : label is "C1DBB623764BA37E2D36331F4263E84D8CE7BD6C0AC207A1C88888CC8CC8C8CC";
    attribute INIT_10 of inst : label is "9262219A0C0B085A084F90A11933951544C218AC3158C5D73133C555ECD3276E";
    attribute INIT_11 of inst : label is "71100F80200E9A1609580C5618AC62E3B9898DE2AAF4901E1E04924924924924";
    attribute INIT_12 of inst : label is "04887012538C3C2442C21610B0858281682B1025310E99799C293A60B09C8AC2";
    attribute INIT_13 of inst : label is "B0BB871A6AC4C006820820820820820C87098169B6E4812009004A02C0168094";
    attribute INIT_14 of inst : label is "0924941666120A47EB0DAE2B1DAAE173FDAE2B5DAAE160C2042130C28EBC3569";
    attribute INIT_15 of inst : label is "E6683799B718E0002A28A4C90B2E42EDB3431456CC08645256AB248F408F40A0";
    attribute INIT_16 of inst : label is "20808A061040C5030820228184103140C20818A061040473227C9328AB36741B";
    attribute INIT_17 of inst : label is "35141841D062B0BAC4104505CB4AA40000D3AA69D5342818020228184103140C";
    attribute INIT_18 of inst : label is "0000000000000000000000800022B1351252484C26A2A24B8ADA40A4FC484895";
    attribute INIT_19 of inst : label is "03C00000C0000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0408004080040800408004080040800000000000FBFFFF000000404080810100";
    attribute INIT_1B of inst : label is "35E62700C4240028000000000000000000000000000004080040800408004080";
    attribute INIT_1C of inst : label is "8E43893263BBF9C0E4924B6362B6992EB6CF039650D7A09764EBB06B43632826";
    attribute INIT_1D of inst : label is "EDB666FACA5C296A1715A9576E176A549750C6756FAED18E48948E49968E4996";
    attribute INIT_1E of inst : label is "1334B3C31985295ACC36858450C6325B6E896DBAC09405A42C212024230ADB8E";
    attribute INIT_1F of inst : label is "1054A2626A4647DB9AA64B00000000000000000000000DA605498A420484FF24";
    attribute INIT_20 of inst : label is "CE5C3878F1C284B364CC284B364CAC438B12CD9338B12CD932B108B93A124864";
    attribute INIT_21 of inst : label is "B475C644558A5194614A2AC14073B226C8AD7A6D460AD37118305414AF4DC471";
    attribute INIT_22 of inst : label is "2946518528AB0501CE889B22B5E935182B49E460E15852BD2711C5228CC89B22";
    attribute INIT_23 of inst : label is "FA595721B0CA84B0C24F21A1A823925F6ECC63A7A0348A32226C8AD1D71D1156";
    attribute INIT_24 of inst : label is "F0CEA72FE5B6E5BFDF2413368327A318CE730C3D6508A4A1227A7A375FB5D5E8";
    attribute INIT_25 of inst : label is "2858311946CC2365591D22E4751B308D9564740582C160B45604802C042C2121";
    attribute INIT_26 of inst : label is "9D0D0D0D0555678B8723AC5C391D46CE2365591922E4651B388D9564650B0623";
    attribute INIT_27 of inst : label is "8A7AE2F66B2D3FFFFEE0000FFFFEE0000CC1CA0054646464640000746474341A";
    attribute INIT_28 of inst : label is "1A8A6A94C5316C53654C5B14D953654C5E7AF59A79EB5736A7AF58A6983A8A3A";
    attribute INIT_29 of inst : label is "B4A52775B335A8B29808172CF2DC266A2496E575E5B237713569515515135695";
    attribute INIT_2A of inst : label is "293AEDD9ED403501AB6ED294BD76ECF6A01E00D5B7694A5EEB666B500F006ADB";
    attribute INIT_2B of inst : label is "7AADCF6A01A00F1B5694A5EFB666B500F4078DAB4A5277DB335A806A0356DDA5";
    attribute INIT_2C of inst : label is "EDD9AD403401AB6ED2949DF6ECD6A01E80D1B5694A4EBB73DA80780346D5A529";
    attribute INIT_2D of inst : label is "A201F00404007ADBB4A52F5DB33DA807ADBB4A5275DB33DA80680356DDA5293B";
    attribute INIT_2E of inst : label is "B848FF70937DFE102A0A0A0A000AAAA00AA0000AA0A0AAA000A0A00AAA0A00A0";
    attribute INIT_2F of inst : label is "0002000000021A10D04C4E0886176D6D7BAE2CB6D9C6319CF0A6D23E4FABB30F";
    attribute INIT_30 of inst : label is "020D800000000000000008000800000100020000002000100000020008000002";
    attribute INIT_31 of inst : label is "06040404000A0E0E0A04000A0E0E0A04000A04060A04000A06000C0400000202";
    attribute INIT_32 of inst : label is "080441042010202208402041010080442EC4108060A0110806082B0080400004";
    attribute INIT_33 of inst : label is "0B0414410884020410110410806082BB10410804020404410804020410177050";
    attribute INIT_34 of inst : label is "CAC964AC964B62100C15D8820840305008840304105762084020410110410806";
    attribute INIT_35 of inst : label is "03C21A02114B4B5A6D6D25253692B69292524ADB5B69A52B4A56B45AD96CAD96";
    attribute INIT_36 of inst : label is "A681A80F407A43C21E10F006803C01A00F006803C21E10F087803C01A00F0068";
    attribute INIT_37 of inst : label is "000000000000000000C0000C0000C00008CE6377C101EE08BB698A27B5C0F407";
    attribute INIT_38 of inst : label is "EF1D947655CF6C7BAD48B6A45A3C00C000180002000000000000000000000000";
    attribute INIT_39 of inst : label is "A6D249B6DB6924924DB6DB6DA4DB486A265364218B162C16D6D6594A5012163C";
    attribute INIT_3A of inst : label is "0080080050200001000016080000683000010480830002000009000420080004";
    attribute INIT_3B of inst : label is "0020020008008088088088008008008008088008088088088088008088008008";
    attribute INIT_3C of inst : label is "8200800000220002200220202002022022022022022022022022002022002002";
    attribute INIT_3D of inst : label is "55555555555555555555555555555555545055555550807C0100000020001040";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555550CA9";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "543622A1B0673B76EDDBB76E993264C993264C993264C9923E7986CCC361DCC1";
    attribute INIT_01 of inst : label is "91138372E1130461C18187869E5C88F13399CCF67B3D9EF37E6FCFF9FF3FE7DC";
    attribute INIT_02 of inst : label is "C6798C13A1301E6FC3ACB4C0621A06838C89031221099C670739CCE733301891";
    attribute INIT_03 of inst : label is "F3058F3180CC06603305982CC1660A301980CC06603305182CCA4233CC666798";
    attribute INIT_04 of inst : label is "166C8473058F3058F3058F3058F01D8C6318C6303058F3058F3058F3058F3058";
    attribute INIT_05 of inst : label is "472265220DB20DB20DB2293329377F83FEFFB5FD83BEA985A7D24D9325A4754C";
    attribute INIT_06 of inst : label is "122932201908832091049984874445B6230C836C83661B187878AAE10E4A5724";
    attribute INIT_07 of inst : label is "301980CC0660318F18CF1E2C8616167210C6DB2926524834D06DB2DA65248249";
    attribute INIT_08 of inst : label is "CC924C3718C16182C23058460B0C602301060208C0418C1660A305180CC06603";
    attribute INIT_09 of inst : label is "0A3050596C32721919832F301A61610D9E398E49949C62B1E12C70E63A4DA436";
    attribute INIT_0A of inst : label is "2C4944E3182CE01CE3324933631B31B523121A4E664C9190C88C187860A0C066";
    attribute INIT_0B of inst : label is "C58E1270B70E700DB613B7938D9C671808F8C806490B125118C6033B87709926";
    attribute INIT_0C of inst : label is "0E953556CB470924B180CEE0C717C6C602398706126405260589320292028738";
    attribute INIT_0D of inst : label is "CCD6365E79B636D98D830E78DC838760D230619CF3404E953E4A3D6767676700";
    attribute INIT_0E of inst : label is "72AA555B2EEAEABA3A3AE0D096DA0017D94379E6DB371B39E364D9CF36DB81B6";
    attribute INIT_0F of inst : label is "2624439C89245B90734B843186C630D8E0412997E6FE60E03777733733733773";
    attribute INIT_10 of inst : label is "8E8B048AC980CC14219AC06606DDCCE339394E4E9C9E32449CB272ABE1349891";
    attribute INIT_11 of inst : label is "9CEFF07FDFF85CE8C800A7274E4F192C24E5B13955F246E268138E38E38E38E3";
    attribute INIT_12 of inst : label is "C169900D28F40C3B60B305982CC168305881C6031C33B1858504C6C251A3E146";
    attribute INIT_13 of inst : label is "06E6D939439F8EFC61861861861861901119301B4D88301180CC0660A3051828";
    attribute INIT_14 of inst : label is "6C924A15BCDB311D467718E667038DD4AB18E627038DD319B187479E50E463E7";
    attribute INIT_15 of inst : label is "3DD8E6F77C9F936B5ADE5234649139304C396F2923312B19055796735B735B6C";
    attribute INIT_16 of inst : label is "96EE737A4B77B9BD25BBDCDE92DDCE6F496EE737A4B773D9BDCF597E606E1C73";
    attribute INIT_17 of inst : label is "8726796699E4F2D3CC150550CA21B6EF6EDB556DAAB7CDE9DBBDCDE92DDCE6F4";
    attribute INIT_18 of inst : label is "FFFFFFFFFFFFFFFFFFFFFF7FFFC4F31B8B7B6C640FE7666C1D0369B62B6C86D8";
    attribute INIT_19 of inst : label is "FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FBF7FFBF7FFBF7FFBF7FFBF7FFBF7FFFFFFFFFFF040000FFFFFFBFBF7F7EFEFF";
    attribute INIT_1B of inst : label is "4152911D06136FD81555541FFFFFFFFFFFFE007FFFFFFBF7FFBF7FFBF7FFBF7F";
    attribute INIT_1C of inst : label is "7B28E1E3C0988C445249067C381C748CEEE51149078881C883244283A7C1A158";
    attribute INIT_1D of inst : label is "324999032120848248420C1890D893109329298190310C7B264B7B27497B274B";
    attribute INIT_1E of inst : label is "44C3617CF45E94B5B9C970DF0F39E936D864DB61182CC1460330589B9C2BE413";
    attribute INIT_1F of inst : label is "431BDB1B27978EBCD5ECDEBFFFFFFFFFFFFFFFFFFFFFF251F0645938C7060598";
    attribute INIT_20 of inst : label is "295983060C132638705932638705D3384C98E1C164C98E1C174CE42D8FC1A190";
    attribute INIT_21 of inst : label is "C305D09305A30C83046182E47736C982E231659C31A32CECC76519462CB3930B";
    attribute INIT_22 of inst : label is "8C320C11860B91DCD9660B88C596F0C28CB7B30D946518B2DECC2F7063660B88";
    attribute INIT_23 of inst : label is "A31C966DC6D899C6CCE16D8D8AC37759D36B5B32DB9DC184982E230C1742CC16";
    attribute INIT_24 of inst : label is "0FA29287136D9095859844CA079058C639CEF1C1902232045B0CC51728D1818F";
    attribute INIT_25 of inst : label is "730364C3C2E131702CC3D8330F0B84C5C0B30F73399CCE6B08C0460B1603305B";
    attribute INIT_26 of inst : label is "B2727272711176606C98730364C3C2E131702CC7D8331F0B84C5C0B31E606C98";
    attribute INIT_27 of inst : label is "9B7ADAC92CAF700000000000000000000FF898001020202020000030303071F7";
    attribute INIT_28 of inst : label is "D2CB889775ED775EB17B5DD7AC5EB17B5B7AC5916DEB96C2C7AC5917BB989B98";
    attribute INIT_29 of inst : label is "421081A30C8347C5CCD27DB32B2398959249129232FC1895B56D5D6D975B56D5";
    attribute INIT_2A of inst : label is "844C58245A36023018910842062C122D1B05182C4A8421034619068D828C1625";
    attribute INIT_2B of inst : label is "4D1820D1B0518084A8421131619068D80CC04254210898B0C8346C0460312210";
    attribute INIT_2C of inst : label is "58245A3602301891084206AC122D1B05182C488421035608346C1460B1221084";
    attribute INIT_2D of inst : label is "5DFE0FFBFFEC06254210818B0C8346C06254210818B0C8346C0460312210840D";
    attribute INIT_2E of inst : label is "18707230ED99ABBC7FF555F5F5F5F5F5F5F5FFF55FF5555FFFF55FF55FF55FF5";
    attribute INIT_2F of inst : label is "FFFDFFFFFFEB05982D35223310EC92909490904924739CF7906D46E5BE8E6CC9";
    attribute INIT_30 of inst : label is "28320000000000AAAAFFF7FFF7FFFFFEFFFDFFFFFFDFFFEFFFFFFDFFF7FFFFFD";
    attribute INIT_31 of inst : label is "0C0E2E2C000E0A082C2C000A0E0C282C000A080A282C000C080E2A2C000A080A";
    attribute INIT_32 of inst : label is "080441042010202208402041010080442644108060A0110806082900806C000E";
    attribute INIT_33 of inst : label is "0B04144108840204101104108060829910410804020404410804020410133050";
    attribute INIT_34 of inst : label is "B1249B1249B122100C14C8820840305008840304105322084020410110410806";
    attribute INIT_35 of inst : label is "60B305886C2626319090D8D8E8686868490921B636C710863188433126DB126D";
    attribute INIT_36 of inst : label is "6C301982CC16603301980CC16603301982CC16603301980CC0660B301980CC06";
    attribute INIT_37 of inst : label is "0000000000000000003FFFF3FFFF00000522912AC6B2225E65C479EC63182CC1";
    attribute INIT_38 of inst : label is "1A204881219633D414124A092543FF3FFFE00000000000000000000000000000";
    attribute INIT_39 of inst : label is "26DB49249B6924DA6DA4DA4DB4DA6F03D109108C366CD9B9090924210FCDC9EB";
    attribute INIT_3A of inst : label is "0880080088200081000830080020683000024D0283000020000A400400004089";
    attribute INIT_3B of inst : label is "0220020008008088008088008088088008008008008088008088088088088008";
    attribute INIT_3C of inst : label is "73DF800000010120002101220002022022002022002022002022022022022002";
    attribute INIT_3D of inst : label is "555555555555555555555555555555555554505055577F83FEFE03C73C71CF5C";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555553E2C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "FC1027E000228000000000000000000000000000000000007E7802AC01514C03";
    attribute INIT_01 of inst : label is "48B90720C0862450A9414503940A48C89148A44221108812A25448891122244C";
    attribute INIT_02 of inst : label is "863888528100B42F82A534C1221200111A44A28911088A228F7BC6C631291541";
    attribute INIT_03 of inst : label is "53008511804C026013049824C126013049824C126093009801880231C4426388";
    attribute INIT_04 of inst : label is "1264045300853008530085300856158C6318C630300853008530085300853008";
    attribute INIT_05 of inst : label is "2492E006001604960016201620100000000137998A2640C72753499325A47215";
    attribute INIT_06 of inst : label is "162016021438096003000B00052C2492E1258125812C09307424AA93491A548D";
    attribute INIT_07 of inst : label is "3001800C0060010A884A9A3A1D15156810024924924924820900000000000000";
    attribute INIT_08 of inst : label is "D800056288C0018002300046000A601300060008C0014C106093049824C12600";
    attribute INIT_09 of inst : label is "083040492A29691491428430405151089E28850B801AD7EBD17C2852292000B6";
    attribute INIT_0A of inst : label is "380022D11820400AD36000152E09609096094EC5264A4B48A48A14226094C106";
    attribute INIT_0B of inst : label is "C7051228F28A2812B21296B14DCA261800D46004000E0008B446001153299002";
    attribute INIT_0C of inst : label is "0C3515529946892491804650A293A646011142853240040204992002000202B5";
    attribute INIT_0D of inst : label is "8E54144820921251A50218225C8183E0C22040B041010C341A0A313333333300";
    attribute INIT_0E of inst : label is "76A8554A66CA82A02022A0D0924AAAB38B5120824A334B60896E5B0416498092";
    attribute INIT_0F of inst : label is "A5122158456C5B50692152170242E0485010424354A220203777773773773733";
    attribute INIT_10 of inst : label is "084B059A41800C1021190AE408018D8363152D4A5A956A404A2028ABA4929448";
    attribute INIT_11 of inst : label is "5A000000003854E8C80896A52D4AB52C0251301455D2C2C27812082082082082";
    attribute INIT_12 of inst : label is "C02980286A7C18336083041820C100304000A6000A2691850485C242709751C2";
    attribute INIT_13 of inst : label is "26A2D833029A9A5451451451451451481708300124A43049820C106013009804";
    attribute INIT_14 of inst : label is "08924E1494D91318026108C261028D500108C261028D531D9345229CD0AC27CD";
    attribute INIT_15 of inst : label is "6118E584741E835AD6556952D44AB490A2152AB4952122140557555600560064";
    attribute INIT_16 of inst : label is "864D4122C326209161931048B0C988245864C4122C326358A15C115D600E1C72";
    attribute INIT_17 of inst : label is "93632B320CAC56415D4005558269124F66495524AA93048B9935048B0C9A8245";
    attribute INIT_18 of inst : label is "000000000000000000000000000C57118939242C0FEE2E2438092B9203258648";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "010AB314060965440AAAAA000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "62A0D183018898C00000023A1434D006A6570000061981A11020020206412100";
    attribute INIT_1D of inst : label is "000000221084420220200A1002D002948100100102201862AC2B62AD2B62AD29";
    attribute INIT_1E of inst : label is "2806203AC28B4A420080684A8E3584800252000B9800C006083000B35A69C000";
    attribute INIT_1F of inst : label is "02194A0A2E1226705F4C9A80000000000000000000002003E852DB3440060B41";
    attribute INIT_20 of inst : label is "294B56AD5AB16225204B16225204F114C58894812C58894813C4502D4D830180";
    attribute INIT_21 of inst : label is "4604C1B6048118862023026036B6DB0240112CB4618165A58264090225969603";
    attribute INIT_22 of inst : label is "046218808C0980DADB2C090044B2D18205969619902408965A580F70C32C0900";
    attribute INIT_23 of inst : label is "3288936C8650DC864E406C8C8AE16748B36B5B2A7B5DC30CB024011813065812";
    attribute INIT_24 of inst : label is "4A96B246480028908B41280E0742F5AD6318C589000220004A06C5126051012E";
    attribute INIT_25 of inst : label is "D6866D86C24311206D82F4360B090C4481B60B68341A0D0E9CC1260116083001";
    attribute INIT_26 of inst : label is "B6D6D6D6D11122D0CDB0D6866D86C24311206D82F4360B090C4481B60AD0CDB0";
    attribute INIT_27 of inst : label is "C93A4A4964A6700000000000000000000008D8003000000000000010101011D5";
    attribute INIT_28 of inst : label is "D25988B3748D3748B1234DD22C48B1234B3A64932CE992C663A44933BB98C998";
    attribute INIT_29 of inst : label is "000001A90D8947A28E0035A22A075441492028068860101595254D24B3595254";
    attribute INIT_2A of inst : label is "000C082C0A36003000900000060416051B0418204A000003521B128D820C1025";
    attribute INIT_2B of inst : label is "0C486251B00180448000003020B028D804C022400000181058146C0060012000";
    attribute INIT_2C of inst : label is "086C0A36083040940000260436051B0018004A0000130218946C006001280000";
    attribute INIT_2D of inst : label is "A000000003EC1025000001A10D8146C1025000001A10D8146C1060812800000C";
    attribute INIT_2E of inst : label is "4820609045B97EB0600AA0A0A0A0A00AA00AA0A0A00AA0A0AA0A00A0A00AA00A";
    attribute INIT_2F of inst : label is "00000000000B0498248566210BA500000034080000E318D6B025C0ADBC0A24C0";
    attribute INIT_30 of inst : label is "0020000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0604040600060200040600060200040600060200040600060402000600020200";
    attribute INIT_32 of inst : label is "080441042010202208402041010080442644108060A011080608290000060006";
    attribute INIT_33 of inst : label is "0B04144108840204101104108060829910410804020404410804020410133050";
    attribute INIT_34 of inst : label is "10124901249122100C14C8820840305008840304105322084020410110410806";
    attribute INIT_35 of inst : label is "6013000848020211000048488024002400801012024500020004221000010000";
    attribute INIT_36 of inst : label is "003041800C006083041820C006003001820C106083041820C106013049824C12";
    attribute INIT_37 of inst : label is "FFFFFFFFFFFFFFFFFFC0000C0000FFFFFC8A450D90226655274C28A5295800C0";
    attribute INIT_38 of inst : label is "0800A002811CA3505C092E04960000C0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "34926D24924DB6934924934D36DB2C13C019000862C58B10000000000FA5A5AA";
    attribute INIT_3A of inst : label is "0880880848200001800002080000683000212000830002000008000021000000";
    attribute INIT_3B of inst : label is "0220220208088008008008088088088088008088008088008088088088088088";
    attribute INIT_3C of inst : label is "0000800000000000000000000002002002002002002022002022022022022022";
    attribute INIT_3D of inst : label is "5555555555555555555555555555555555545050555000000001041800020021";
    attribute INIT_3E of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_3F of inst : label is "5555555555555555555555555555555555555555555555555555555555553E7A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
