-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "54292AA049326940A502940A502940A502940A502940A5007E732429B203E993";
    attribute INIT_01 of inst : label is "089B026254A2AE108B0803128C0B448AA5128944A251283666CCD99B33666CED";
    attribute INIT_02 of inst : label is "9679A95BD064CC6F8A80FDC8D732815B0B00300115AC89A25DEF6667116A3010";
    attribute INIT_03 of inst : label is "C72AEC03953CABE54F2AF953CABE55F2AF913C8BE44F227D3A959733CD4F679A";
    attribute INIT_04 of inst : label is "306C14072AEC72A6C72AEC72A6C4018CE338CE3272A6C72AEC72A6C72AEC72A6";
    attribute INIT_05 of inst : label is "A5508B3651B211FA11B212B212B22B56359FB06185CCBF0DFF1E79F3F43E51E1";
    attribute INIT_06 of inst : label is "EC51FA166C214BA10B28590859F4A599A53E863E863EA1F48A9B2FF0AD016F80";
    attribute INIT_07 of inst : label is "6F0FF873C2BF5CF2F57573054AAE020928A11302CBB5DE4B2ED7790CBB1DE432";
    attribute INIT_08 of inst : label is "9F4FDE8F83D3F4BC7FEA9E55F2E7C77CB9645B9C5B385FC29F5DFAEF837E89E4";
    attribute INIT_09 of inst : label is "19A5A99B295AA55DA82458FA69A69249162C5014094BD1B7A760E4ED5C9D85E8";
    attribute INIT_0A of inst : label is "6CCAE5825A012A20408562F5C9EBDE5CFAB60B0260256400108C7AF40213980A";
    attribute INIT_0B of inst : label is "9678973FD5A248A096591525DEBD36044D2D96410977AB4A012B264B7EB7E813";
    attribute INIT_0C of inst : label is "7A555D373AE79AEE44913038AAEB3D3A41490110C95A16934C9AE64F2D64183D";
    attribute INIT_0D of inst : label is "B4856B8E7CEBCF5C00288523264D9F9C280251145E357A6E79C7AFAD8D8FFEB5";
    attribute INIT_0E of inst : label is "5F5574DBFEBF85210AE666F9FA22CEB765AE1D79EC278A84D53D116F3F275E75";
    attribute INIT_0F of inst : label is "018C863FE303B94402C02212F00F4F15FEB9133A51FA4A3F648639D324F7A37A";
    attribute INIT_10 of inst : label is "DA3E776A924924924924924BCAAD79FC8FF4FB98CBAC5089225170C42188462F";
    attribute INIT_11 of inst : label is "58DA7E2761FFF9D5F69357CA6B56359EDC3BFA1814310862118BE40633818FF8";
    attribute INIT_12 of inst : label is "6BDC8BF4CF26F933C9BF47F22CE6A6AE5D237CF813C1BE44F2651CBD152795B2";
    attribute INIT_13 of inst : label is "6C35CE6E5FA5FF53117FF585513E6D4D61C5EE164964964964964B5559FC8FDE";
    attribute INIT_14 of inst : label is "D8E08920FF1050FB30FB3D27FFFFD80E79C1CBFDB9D65DB9D064B07FD6DDA9D0";
    attribute INIT_15 of inst : label is "78EF31A300C0057A4FCF586C44B8B11DE7BCCE7301625EB5C0AD2782AD00B001";
    attribute INIT_16 of inst : label is "76897E3C7E897E1E3B049F0F1F824F878EC127C3C7E897E1E3B44BF0F1FA25F8";
    attribute INIT_17 of inst : label is "ED6F5FB54A5BACEF4DACFDAB7D5AC6F56FB5DEDAB57D7FB7FE371CFDDFFECFFF";
    attribute INIT_18 of inst : label is "4D6224588856F61F747220F414BADDDCC06D4BD2B5A528CBEDB72B13FADBC93F";
    attribute INIT_19 of inst : label is "A02A0AA02A06A02A06A06A0657403554EAE510A76BB2E5516FD51524575289F5";
    attribute INIT_1A of inst : label is "A81A81A81A80A82A80A81A80A81A81A81A81AA02A02A06A02A06A06A06A06A06";
    attribute INIT_1B of inst : label is "B5621B1FFF9749BD8492174BBF95FEFB64B3DF6DB6E11FA81A80A81A81A81A81";
    attribute INIT_1C of inst : label is "022759AE44C44AE2B2072BAE440E1CAD6A2EEAEB7594FF6AB5AD9257AD4C8EAE";
    attribute INIT_1D of inst : label is "8E3472AD9518EDB28EB1C33A8E4BA382305F6CAB3757AB6DDB8BD59526569A19";
    attribute INIT_1E of inst : label is "0000020000400002060001D2F50E6CA2248525CEE5B22E75A1447395EAF578E7";
    attribute INIT_1F of inst : label is "000001E1F999554001D4B2555560020220200202000048000284000000028400";
    attribute INIT_20 of inst : label is "E0100E8100E63B19676F0C4142D50066E235C073A8DC00AAA001C00AAA000000";
    attribute INIT_21 of inst : label is "A5040400440000044063B19620000E8080E0080E8000E0000E8000E0100E8100";
    attribute INIT_22 of inst : label is "909BAD0067BFFF7F7F7EFFFF6E4151111040475840B2D9750AAAAAAA5555556A";
    attribute INIT_23 of inst : label is "A2BA32D2DD34DE93D6E9A43134A5B4B70A7791CF3C71C71CF3CF1E63484D2020";
    attribute INIT_24 of inst : label is "496D8E1CA50070E591282838183831292939193924A9249249000000000842EB";
    attribute INIT_25 of inst : label is "40B748903917C99F06F86783BB521C19004923833E39F1CF8E7C7BE3DF1EF0F6";
    attribute INIT_26 of inst : label is "DF10D08421084A722ADE12D00000004A62A8DF10D08421084A72AAEABFAAEAEE";
    attribute INIT_27 of inst : label is "21084A622ADE12D00000004A72A8DF10D08421084A72AADE10D00000004A7228";
    attribute INIT_28 of inst : label is "2ADE52D00000004A72A8DF12D00000004A72AADE12D00000004A7228DF12D084";
    attribute INIT_29 of inst : label is "37E9BF0DF87FC3FE1FF0FF87FC33E1BE52D00000004A6228DF52D00000004A72";
    attribute INIT_2A of inst : label is "E9A0E4CF26F937E99E4EFA67937C99F4DF27FD37C99E4CF26FC3FE1DF0DF86FC";
    attribute INIT_2B of inst : label is "00048924916EDB6DD80000006EFA79D80820804EDB6DD40000007EDFEDFD6937";
    attribute INIT_2C of inst : label is "304084059BAD58D67B00000007EDFEDF40000016E9A69D80820006EFB7DD8000";
    attribute INIT_2D of inst : label is "55C05921214AC02D15D5CA592120557116480812B00B45758AE9A313AD600000";
    attribute INIT_2E of inst : label is "E65042D1CE9CB7E333EEFB9B014B67BA72DD8DCDBB5200D91351042DCB624045";
    attribute INIT_2F of inst : label is "9B014B67BA72DD8DCDBBEE65042D1CE9CB7E333EEFB9B014B67BA72DD8DCDBBE";
    attribute INIT_30 of inst : label is "719B6372AB8301CB570609820571AB8715C55C38AE2A05D349B8CE338CD722FB";
    attribute INIT_31 of inst : label is "5EF1978E4E3978E4E39618E6B40B062AE403C1EC19F07B8CF83DC67C1EE33E0F";
    attribute INIT_32 of inst : label is "C143E8A2034D02B5332CED4694400A0140200504A24333A85817F8026116AE8E";
    attribute INIT_33 of inst : label is "BF8FC56BF28AA94658C0000258922589225D45CF690BD29282118AD000003A93";
    attribute INIT_34 of inst : label is "A187A94CCAA3198840E9C74E621030EAAA8000001F6CDB55D1655FC47BB97942";
    attribute INIT_35 of inst : label is "0E6B4087FFFFFFE5151DBA7C2ADE45181856A0AFC2EA6B5398A8AAEFBD7B5150";
    attribute INIT_36 of inst : label is "E633BDF2ABAB1E5ABAB163A0CE3575E371575E3E5C101F4C9801C1A6887C4162";
    attribute INIT_37 of inst : label is "5CEB3A576664666451E27319F1398CF89CC67C4E633E27319F1398CF89CC67C4";
    attribute INIT_38 of inst : label is "CB72D788BF5124BA96D6B416C9015C9095CD7B2406484C07901FA8925D4B5090";
    attribute INIT_39 of inst : label is "EAAB4AFCA2AF98BF552CBB96D6B404C9095C9015CD7B2426480C17901FAA965D";
    attribute INIT_3A of inst : label is "6362430000065A5C297696896363C9C3D955D19974FB79C8621881BF0091E95C";
    attribute INIT_3B of inst : label is "4544111911911911B30000000000191E1E1E0E0014AFEAF4CF1D31ADDBB76E43";
    attribute INIT_3C of inst : label is "FDF7D77755D77DFF777D75D5D7DD500040400404001440444445150111111044";
    attribute INIT_3D of inst : label is "FA92335AB1ACFDCD0326F4B77240893D2DF34A9F2429FFFFFFFE0000001FDD7D";
    attribute INIT_3E of inst : label is "2C0E5CF7F142DA31A5CF1C0530B1C39110AEEBF0761CB09A350BDDEAC54C94B0";
    attribute INIT_3F of inst : label is "D60F0434030600489B447BB79FFA382509C5910075B5155DA3274C0E28B4A1BB";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "03F0E01E96662CCBB32ECCBB32ECCBB32ECCBB32ECCBB32CC0834C91864F9187";
    attribute INIT_01 of inst : label is "2CF32666DAC6F65DBD6B7727FCDA3AE66E3F1B8FC6E3F128CD18A334628CD19C";
    attribute INIT_02 of inst : label is "077D90551A61BC80178276170086AA333A6672448A9198560779CEDEFB0E7279";
    attribute INIT_03 of inst : label is "F8500FB82841400A005082841400A105082841400A005086843800BBEC8477D9";
    attribute INIT_04 of inst : label is "11AB2E78508F8508F8500F8500FD9FC0701C07008508F8500F8500F8508F8508";
    attribute INIT_05 of inst : label is "18F271A485004548450047004700731029BCB2ED8FF89D40E820820C089B74F3";
    attribute INIT_06 of inst : label is "36852440049312444242122212D8016F6C58111B111B08DB17833FF4404607A7";
    attribute INIT_07 of inst : label is "825892CC9605B925C05F084AC1E8A4A70DA87EB4104A21B0D369A24104A21B0D";
    attribute INIT_08 of inst : label is "01A80340B0681242C03724F927813CC97009D2C1D242E41760B305802C03720B";
    attribute INIT_09 of inst : label is "246C1CD258C7E3D2BD62D10C96C9EDB634E9395ED7B42800542C1A04C3509615";
    attribute INIT_0A of inst : label is "097FED1A11270FB28913640A803421A2050878E944E1D67B224C8D00CF48C25E";
    attribute INIT_0B of inst : label is "B1A984E02A0604DB021248E16140164EC7C88492385850036B18DBD91B1122C9";
    attribute INIT_0C of inst : label is "349577C80BFBEEB0B00B02796E92C2E024D8926B18C76E30B5849EC0D8592CEB";
    attribute INIT_0D of inst : label is "F3D24F34B592102CC98D369618F0C424993D1A7BE1DE3496204B33311111555E";
    attribute INIT_0E of inst : label is "AC55DF22FEFFB3B3B3624292D5F7B3C3C93CF2421450BCCA1685A78A5A0C9082";
    attribute INIT_0F of inst : label is "839FD67FEDCE2022CC8891B182240F23F8703102C448788DAC577FF56C394C34";
    attribute INIT_10 of inst : label is "6080F01F0830830830830832855D1601605A80424FE63250343301C8A3990E63";
    attribute INIT_11 of inst : label is "02049E465C4E840101B00416331029BC4C94B55C787228E643980E0E7C359FFB";
    attribute INIT_12 of inst : label is "9E23600F805D06C03721B005884B41C780495113A09404E02741A3529A606856";
    attribute INIT_13 of inst : label is "95481089C6C0208C2C400879ECC4F2359397FC8820C30820C30822AB04016071";
    attribute INIT_14 of inst : label is "82111D91FF59227002700A43FFFF051CFE929BFAD3695AD36995C8FF695AC369";
    attribute INIT_15 of inst : label is "5A9079E449E42F4AE88020A59A411666EC5D08620B413A72CB9CB30ECC85A1B3";
    attribute INIT_16 of inst : label is "58F64CAD48F64C56A07B262B503D9315A91EC98AD48760C56A03B062B501D831";
    attribute INIT_17 of inst : label is "2FAE07BF14AA01F895B20CB568AA8BE6AD557D501F75DEFA27CBD2B12DFF92FF";
    attribute INIT_18 of inst : label is "DB83EDE0C4B0C4B1A6431E2EB9A411199C0B6080200802A26F57FC280036A060";
    attribute INIT_19 of inst : label is "D75D75D75D75D74D74D74D71181B78FF8A878A7B5C74863C5BEE3FF8CA63C4CA";
    attribute INIT_1A of inst : label is "75C75C35D35D75D75D75D75D35D35D75C75C0D70D75D75D74D74D75D71D70D74";
    attribute INIT_1B of inst : label is "06CB7D029A33A0560F40B3A2541AEB6CAA256D925F5CB375D75C75D35C35C35C";
    attribute INIT_1C of inst : label is "C914FE1812DDF03967B1C01892E343FCB80C8DB04FE6D66C06F03C91019DE8DB";
    attribute INIT_1D of inst : label is "41300B0899981F130169AC0C010BC0564AE331FC62F95CE4317CAE7FF9C944BB";
    attribute INIT_1E of inst : label is "FC007E42423C007E02020110EC956125024A469A65121578900680590D86C012";
    attribute INIT_1F of inst : label is "000001FE1554000001E1612666610A50A508407E4A4A04003FA323FC003FA323";
    attribute INIT_20 of inst : label is "E8180E0100EC319C31E60800874A0054D001A41B6000010CC0000010CC000000";
    attribute INIT_21 of inst : label is "CC00000404000004048319C348080E0080E0000E8080E8000E0000E0180E8100";
    attribute INIT_22 of inst : label is "A53F7FD2AE880888888019111900EBEBE940434D74C35669A19999999999998C";
    attribute INIT_23 of inst : label is "55F0898083E04C09ADDBFB7B7F83406967CBC30D34D30C30C30D32CE5C7D61F3";
    attribute INIT_24 of inst : label is "979671B917978DC83508282808283509292909292504924924ADB6DB6DB5AD1C";
    attribute INIT_25 of inst : label is "FF6FEFA952A49404A225406AD7F7E356F7F7DC6AC1760BB05D82E41720B90DC9";
    attribute INIT_26 of inst : label is "1DBDF9CA729FBF0F161DBDF9CA729FBF0F961CBDF94E5397BF0F142ABFFFBC7A";
    attribute INIT_27 of inst : label is "729FBF0F161DBDF9CA729FBF0F961CBFF94E5397BF0F141CBDF94E5397BF0F94";
    attribute INIT_28 of inst : label is "141CBDF94E5397BF0F941CBDF94E5397BF0F141CBDF94E5397BF0F941DBDF9CA";
    attribute INIT_29 of inst : label is "E89764FA27C12E09724B825C92E09F0DBDF94E5397BF0F961CBDF94E5397BF0F";
    attribute INIT_2A of inst : label is "5BFF5B925C96E4B704B82DD12E09725B925C96ECB704B82DC13E89744BA25D92";
    attribute INIT_2B of inst : label is "244EADB6DDA249244A209044A2CB044A2CB2C4E249245E2402408240240A968A";
    attribute INIT_2C of inst : label is "79DBDEDE7DCC40A6F60240240E240240E249245A2CB2C4A2CB044A209044A249";
    attribute INIT_2D of inst : label is "FDD2A85E55BCC5BE78EE6CA85B54BE75AA16D52F316F9E3E5C8D717C9AE4924A";
    attribute INIT_2E of inst : label is "81AAAB7C78D5E18E85080204AAEDD16357863B1420A2A3003636AAB64DA094A6";
    attribute INIT_2F of inst : label is "04AAEDD16357863B14200813ABB7458D5E10EC5880206EAADF1E357843A16200";
    attribute INIT_30 of inst : label is "970604E717DA699E2FB4D93416671FDE6D98FEF36CDBB6AA7F3B80E0B81E4F82";
    attribute INIT_31 of inst : label is "B596B8B6E2DBCB6F2DB8238ADA53E7FBC8FE8853F02214B8110A5C08852E0442";
    attribute INIT_32 of inst : label is "09D7BD655ADFDF6EAAC58F2FA0C89913626C4C8FC791760B18C5B9A68C39DD78";
    attribute INIT_33 of inst : label is "66A18FD1FD9DD811338924AEE3B8EF3BCEE5CF20DC3018DFDFB39F824929E788";
    attribute INIT_34 of inst : label is "D75C00BB8D607714981508A1C526EB99999C243A4A80212022B1AE0A73323ECF";
    attribute INIT_35 of inst : label is "F8AD851C22222256622340024C848A2CA4E0CC7027207C6E713115530A021A6B";
    attribute INIT_36 of inst : label is "8AE0636717F26CF17F264E256CE3FECD663FECCFD9DDAAA9773FF377DC88AE9D";
    attribute INIT_37 of inst : label is "E02C0DFC8D8D8F8FEF45C57022E2B811715C08B8AE045C57022E2B811715C08B";
    attribute INIT_38 of inst : label is "6D9B63C5873AD5E0DB05E29B02DAF02DAF38B60B6816D429D4839D6AF06D9922";
    attribute INIT_39 of inst : label is "C7FFB47F6773C5873ED5E0DB05E28902F2F0252F38B60BC8129439D4839F6AF0";
    attribute INIT_3A of inst : label is "FED7D7EDB6DFA3F69577EA8817D6829C2A3BBBFE3F6D5F136631CA1F5ADB36F0";
    attribute INIT_3B of inst : label is "1051190999998889B3800000000050E62AAA96000F92F88774947FF76ADDABDF";
    attribute INIT_3C of inst : label is "55FD557D77F55FDD7D557F55FD5FCCC844CCC44C8CC450455054114401544055";
    attribute INIT_3D of inst : label is "4E055798814DE25FCB82606897F2E0981A17D9F17D9F1FFFFFFE00000017F57F";
    attribute INIT_3E of inst : label is "4074EB0A1A3C3C8550EDD6C0E70F8EFD74BFC6BAD394E69A9C094870E701AD6B";
    attribute INIT_3F of inst : label is "8822A7CC850A2C1061358CFE294B426F56FC8F26D8F939213E3E1404E2AC98AE";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "55E6CAAE2745BB74EDD3B74EDD3B74EDD3B74EDD3B74EDD07CC90CE4A6729C86";
    attribute INIT_01 of inst : label is "9BAA054093A4A8716ADBC21508548AF135D2E976BB5D2E5B23646CAD95B23651";
    attribute INIT_02 of inst : label is "C451384B0321E8628501B7F60EF4381A14DDA7BB752D56B58A50A8A522F26893";
    attribute INIT_03 of inst : label is "A7D4AA23E81F50FA07D4BE85F52EA07D0BEA5F42FA97543A84A80EA289E24513";
    attribute INIT_04 of inst : label is "001D0A67D4AA7D4AA7D4AA7D4AA1181C0701C070FD42A7D42A7D42A7D4AA7D4A";
    attribute INIT_05 of inst : label is "A23113A91500154815001548170012E0A15E20AD26FA0AE1A30EBF76ED9A7051";
    attribute INIT_06 of inst : label is "48954810B0C552C1D48EA40A80E32B249503055207522A01856A4AA528534569";
    attribute INIT_07 of inst : label is "85F9AFC9566ABB55D264EF45B0D03032C10876916DB09241B6CA4D94920DB612";
    attribute INIT_08 of inst : label is "2FA05F5093EA133FC1D70BBA5DD2FED7E4E8A7D8A7FFE5FF0EF17783AC5D72EB";
    attribute INIT_09 of inst : label is "732B0DD496B55AA5945AA0FB4D26B259293FDEE33DA7EA57D4A4FA149F4299D4";
    attribute INIT_0A of inst : label is "5B548A00CED2D2C9DC9842EB05D70EB07588D74C3A5A5919932875C260677A15";
    attribute INIT_0B of inst : label is "2C556EDBAE05B810B600775BBF60F58AB225849DD6EFDC3842D66D2B493493B3";
    attribute INIT_0C of inst : label is "6CC01F6D160C35DFB072D386651F7AE1E7569D11D6B41A2D4D6BD8B776ED385A";
    attribute INIT_0D of inst : label is "E918F1CF4AC9657A0CF3C3F01C39D144C98FE78EFECB6CEF08B1999BBBBAAA8B";
    attribute INIT_0E of inst : label is "AE007DB7D53549C9C0E1003D257D3976CFC7192CB8FF471FE3FA78F7A4164B27";
    attribute INIT_0F of inst : label is "0D6F05B54E9843DDB8776E2D6DC37A681F84AC4955242AA48B075CEC4B2DA83A";
    attribute INIT_10 of inst : label is "ABBA955D144105144105144609A8505F72AEA77A424698CC922AC6B4AD613588";
    attribute INIT_11 of inst : label is "BAC8E04158313014492C513592E0A15F1096B7444DAC2B584D62A8B5BEA16D53";
    attribute INIT_12 of inst : label is "6B3D42EB975C3EC1F62FB97D80EB536C110B05AEE9774BBB5D903D70025BAE05";
    attribute INIT_13 of inst : label is "EA715A9DB719CAD13913CDCB3BBEC354ED690B145104104145145635425F70DB";
    attribute INIT_14 of inst : label is "BBD12E29AA6180D480D000419249950B21F15553BBDEABBBDCEA70AADEABABDC";
    attribute INIT_15 of inst : label is "3665A0E188E00A80F805508F72A13DC1EA3DA94B0286DBACF6EB631BAB01436D";
    attribute INIT_16 of inst : label is "6CBD1A9B3ABD1A4D9D1EAD26CC8F56936747AB49B32BD1A4D995E8D26CEAF469";
    attribute INIT_17 of inst : label is "A2A0D88A96C86D04DC39B73D1DE9DD33A3D3A7423FD7FC95E56F4A7BF754FBAA";
    attribute INIT_18 of inst : label is "4D71945C47EF3A8AAF5111D0AC57EE944A240635AD635819A3D0D436C6D8C847";
    attribute INIT_19 of inst : label is "BE1BE0BE0BE4BE1BE5BE5BE4E9126C2808A30622B47BA233B4EB4A0110518706";
    attribute INIT_1A of inst : label is "2F92F96F96F86F82F82F92F86F96F92F92F92BE1BE0BE4BE1BE5BE4BE4BE5BE5";
    attribute INIT_1B of inst : label is "2DA8DC2196396E7EF2DCB9687CC7075DC684EBBFEBA6396F92F92F96F96F96F9";
    attribute INIT_1C of inst : label is "22A0A12095910E84D4203A2015AB5651055003420A110A83A05336E6E8150034";
    attribute INIT_1D of inst : label is "527493A75D3924EB9254AB435218A489B29CE65322E7539C9173B9CA0314DCAA";
    attribute INIT_1E of inst : label is "FC003E42423C007E02020107490B97E1FC693F490CEE76141536B49D6EB71922";
    attribute INIT_1F of inst : label is "0000000019995540005354C787A10A50A508403E4A4A04001EA323FC001EA323";
    attribute INIT_20 of inst : label is "F0180F0180F6658EB9D10C00439C00585040A0814100000F00000000F0000000";
    attribute INIT_21 of inst : label is "0304040044000004402658EB18180F8100F8180F0100F0180F0100F8100F0100";
    attribute INIT_22 of inst : label is "99DABD98A0955DD55DDD444CCC4014015420945424020814507878781E1E1E0F";
    attribute INIT_23 of inst : label is "4D92A991B364648CA6C9B3ADA4A32465B6C5BA68A28A69A69A68A23444951253";
    attribute INIT_24 of inst : label is "01A43EE021A1F703BF2A0A1A3A1A1F2A0A1B3A1A065B6DB6DB3B6DB6DB39CE93";
    attribute INIT_25 of inst : label is "4D352918EEC5760AB055C3BE08687DF040690FBE1DC0EE87743BA1DD0EE07701";
    attribute INIT_26 of inst : label is "22B99C6339C633FC1822BB9C6339C633EC9822B99C6738C633EC982ABFFF96DB";
    attribute INIT_27 of inst : label is "18CE33EC1A23B99CE718CE33EC9A23BB9CE319CE33EC9A23B99CE319CE33FC1A";
    attribute INIT_28 of inst : label is "1822B99C6738C633EC9822B99C6738C633FC9822B99C6738C633FC1823B99CE7";
    attribute INIT_29 of inst : label is "C95E6AF25792AC95E4AF2559AACD5E42B99C6738C633EC1822B99C6738C633EC";
    attribute INIT_2A of inst : label is "C9B4AB35D92ACD766AB35D9AEC9766BB25592EC9564BB35592BC9566AB25792B";
    attribute INIT_2B of inst : label is "4916ADB6DDC892491488241148834D148D34D16892491C090091C09009024403";
    attribute INIT_2C of inst : label is "B1A46723294B82857E40900904090091E892491C8D34D148834D148824114892";
    attribute INIT_2D of inst : label is "B116E5EF78FA91BFB5B7A7E5EA79ED44B97F9E7EA46FED691FBB60A8D68F6DB7";
    attribute INIT_2E of inst : label is "B3B7F1BBEBB14BA9DFBBAECC9FC6EFAEC52EA77EEEFB4D72DB7A7E1B86CBDEE3";
    attribute INIT_2F of inst : label is "CEDF86CF2EC52CA67CEEBB337F1B3CBB14B29DFBBAECC9F86EFAEC52CA67EEEB";
    attribute INIT_30 of inst : label is "36CD2775BAF765D575EEC3B0BC7EB2F365FD979B06C99CF3D68366D9B645952E";
    attribute INIT_31 of inst : label is "E9192CCAA32A8CAB32A97B4EECD8D1B0B0E574256CDD09B66E84DB37426D9BA1";
    attribute INIT_32 of inst : label is "CCE7D934CA4D9334376E486CCA0E43C8390720E66F479B891245A4A5C42D9BB4";
    attribute INIT_33 of inst : label is "C60C4ABB5C1F965534B6DB70B4290A42D0A777EF92DBB6749CAD616DB6DEFD6B";
    attribute INIT_34 of inst : label is "7492A1F74F876E9CD19B4CDBA734DB4787968F68EFB1743737E4EF1F4AAD6F0C";
    attribute INIT_35 of inst : label is "B4EECDDAEEEEEE633332D21EF1EFDF78FAB270FBE58E46394B9999F9DF638B33";
    attribute INIT_36 of inst : label is "4ED95275BAFF6EABAFF6EC8D8FD65F6F7F65F6EB4D88B3CDEE9CE3C515D7619B";
    attribute INIT_37 of inst : label is "F45916A87C6C7E7ECDBBA76CDDD3B66EE9DB3774ED9BBA76CDDD3B66EE9DB377";
    attribute INIT_38 of inst : label is "4FD1B001B167C7461F85420DAFF3A2F53A37FCBFCD7A9C3C0498B3E3A34FD3F4";
    attribute INIT_39 of inst : label is "2515F2D707E001B163C7461F85421FAF7BA2F7BA37FCBDED7BDC2C0498B1E3A3";
    attribute INIT_3A of inst : label is "6E676632492620A2820A28A0808AA2082CB362EF6D23BE9A84290FB5890A9AA0";
    attribute INIT_3B of inst : label is "EBAEAA23223323220180000000001088CCF712001275C5D4CBCE631CB97AF646";
    attribute INIT_3C of inst : label is "8A2A082A88A88A002A8A2808A08A15D91995D19995FAABAFAAFBEBFABEBFABAF";
    attribute INIT_3D of inst : label is "1174B697050AF1E89E2324647A2788C9191A6DB1A6DB00000001FFFFFFE8A88A";
    attribute INIT_3E of inst : label is "2A0995C5D5C35383289424B1201880A3098712892B2C5F34020184809CBD4C52";
    attribute INIT_3F of inst : label is "D041433272E7C38F24ACE23DBFBD59D227CE430C33A3C383C7C7804609AEB50A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "BC5325E299DC64C993264C99326DDBB76EDDBB76E4C99324F80B28B594586D93";
    attribute INIT_01 of inst : label is "664E20C40A70694A1A352A3828A135E6582C160B0D86C3542A8550AA554AA954";
    attribute INIT_02 of inst : label is "10820154CB6488A597B3FC0484A6A33E3176EEEDDA03314848021088660E2665";
    attribute INIT_03 of inst : label is "081A90880D407A03D01A80F407A03C01A80F407A03501E00F5A814A4900B4920";
    attribute INIT_04 of inst : label is "11092D481A9081A9081A9081A90D522A8AA288A201A9881A9881A9881A9881A9";
    attribute INIT_05 of inst : label is "5DA26F8074027426742675027502441F004083DC1B33E447A324D3AF4D9AFF23";
    attribute INIT_06 of inst : label is "92F502701AB3C027427A013A8109E976DF009D099D00EA061716BAAED7EEBD37";
    attribute INIT_07 of inst : label is "401680B405802C0160024A4A09C42C2E25A98924B6DB2CB6CB24B2C92CB6CB64";
    attribute INIT_08 of inst : label is "803C0078580D0AC0B005802C01600B0058488A508A409404A02D01600B004802";
    attribute INIT_09 of inst : label is "A6509FC02108068A4085890D9659E9A662E96B5EF6B40F401E9603D2C06A5606";
    attribute INIT_0A of inst : label is "09C49894836E2E366B57C4024005A0240163504B0DC5C6CD6AF88169585A5240";
    attribute INIT_0B of inst : label is "438714840B0C505A2E015DC520585C798AC3805771481611462199BF09F09ADF";
    attribute INIT_0C of inst : label is "A2AA92082959609025263AC31442409095F1D64231094042B2149308C349AC8C";
    attribute INIT_0D of inst : label is "22124D36DADB4D08E94D32426A13C11295249A685574A2AE2159111111114034";
    attribute INIT_0E of inst : label is "1CAA482054D532B2BAEB4E1B62A0528A2934DB69944934C92249A6936E76DA60";
    attribute INIT_0F of inst : label is "73133C555ECD3276EC1DBB621760BA37E2D36331F4263E84D8CE7BD6C0AC207A";
    attribute INIT_10 of inst : label is "A4A4F2F02492492492492493114CD0E0580252527C847141504C218AC3158C5D";
    attribute INIT_11 of inst : label is "53A65E670A0E980C2722309C441F004174D4B44AC062B0C563175DCC4D6F1557";
    attribute INIT_12 of inst : label is "B9207802401680B404A02501625C0495E30F0900900480240120A05A0AC40B4C";
    attribute INIT_13 of inst : label is "BA58B489084D34ABAF0D5A752EE5C6AAB53421A08208208208208329C2E05A6D";
    attribute INIT_14 of inst : label is "12991595AAD963D023D0280249250599A40215FAD36BAAD76ABA5CFF6BAAD76A";
    attribute INIT_15 of inst : label is "0808E644F9262A2ACD9D26F99A4DE66DC638000A8A2B7242DB90BB6CD0C515B7";
    attribute INIT_16 of inst : label is "685234040C52348206291A4101148D20818A469040452348206291A4101148D2";
    attribute INIT_17 of inst : label is "55549755B48549F892912A56A83483A0D56975AA8A28AB9685490011A754D3AA";
    attribute INIT_18 of inst : label is "000000000020A50402040000A02809000090400420080004156A6A24A490984D";
    attribute INIT_19 of inst : label is "104104104100104100100100228960D32008425849100000904034D8CA040004";
    attribute INIT_1A of inst : label is "0400400400410410410400410400400400400104104100104100100100100100";
    attribute INIT_1B of inst : label is "01494F904164505208A0ED505208400005042080080CA4040041041040040040";
    attribute INIT_1C of inst : label is "C19F571A128CB418A592D01A12A549AC9029C690F572824503A1840B409D7C69";
    attribute INIT_1D of inst : label is "00000000000000000000000000400016428092501002009208010034D8CAA0BA";
    attribute INIT_1E of inst : label is "0000000000000000000001F00000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "000001FFFFFFFFFFFE0000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "08100081000000000001FFFFF800000202040408081C01FFE001C01FFFFFFFFE";
    attribute INIT_21 of inst : label is "0040004400044004400000000810008100081000810008100081000810008100";
    attribute INIT_22 of inst : label is "2D6792728F919999911111199110000000061040820060040000000000000000";
    attribute INIT_23 of inst : label is "BA7E84F4A99D0BA55992DA4249E07C0EDB2C612010012482480410DE1B286CAB";
    attribute INIT_24 of inst : label is "B6B6D035129281A13606061406061607071407071164B6D924E4B6D924A76BEE";
    attribute INIT_25 of inst : label is "B2CDA56940F007807D03E00F0DADA06A24A4940D007803501A00D406803D01A1";
    attribute INIT_26 of inst : label is "C887294AD6B5AD4924C885394AD6B5AD4924C887394AD6B5AD4924FFD57FE954";
    attribute INIT_27 of inst : label is "D6B5AD49A4C885394AD6B5AD4924C885394AD6B5AD4924C885294AD6B5AD4924";
    attribute INIT_28 of inst : label is "A4C885394AD6B5AD49A4C885394AD6B5AD49A4C885394AD6B5AD49A4C885394A";
    attribute INIT_29 of inst : label is "B005802D01600B405A02D01680B005A885394AD6B5AD49A4C885394AD6B5AD49";
    attribute INIT_2A of inst : label is "12DB02D01600B405A02C01600B005802D01600B005A02C01680B005A02C01600";
    attribute INIT_2B of inst : label is "000000000800000000000000000000000000000000000000000000000000B4DB";
    attribute INIT_2C of inst : label is "FDC9DADF87107C01000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "5A0AB080528F25D2DA9B983094529682AC2014A3C974B6A794449382C32496D8";
    attribute INIT_2E of inst : label is "ECD898671C5C1C1178EDF3B362619C71707045E3B5A0C3E826A488879801009A";
    attribute INIT_2F of inst : label is "912221BCF1307044E397CE458986F3C5C1C1178EDF3B362619C71707045E3B7C";
    attribute INIT_30 of inst : label is "8C10D4A34E4AC88E9C95996652234E4ACC8A7256659D529A2466098260B4F071";
    attribute INIT_31 of inst : label is "823483A50E947A51E947220949567CE69AB89B924326646093323049991824CC";
    attribute INIT_32 of inst : label is "0DBA24E3AC96CCCF4C91A2F12CAC9596B6D6DAD9148E672D2B49BA9A94C84260";
    attribute INIT_33 of inst : label is "F79FBD754B5441D099896DA50942D1B46D1CCBB006354F49A9C21C325B69F01C";
    attribute INIT_34 of inst : label is "78A24AA21646441AD9A4CD3706B78600000000070AFC26EBA292AAAA9446A5AB";
    attribute INIT_35 of inst : label is "6094B570000000433334761004E46A3ABCA507D59519922109991111CAAAEA35";
    attribute INIT_36 of inst : label is "098204234E5AE474E5AE5F95C469CB5F229CB5ECCBEABA29C19393F84089B426";
    attribute INIT_37 of inst : label is "A0A5390281818383634D04C1268260934130C9A09864D04C326826093413049A";
    attribute INIT_38 of inst : label is "92A589F37E59B819254812618402084020A09610082013E39BBF2CDC0CD2B58C";
    attribute INIT_39 of inst : label is "DAEACD52D51DFB7E59B819A54812618402084020A09610082013E39BBF2CDC0C";
    attribute INIT_3A of inst : label is "949494A496DCAA40A882222888A2208A02C84BDCA77ABC139AD6B254CF57500A";
    attribute INIT_3B of inst : label is "DD7DE323322222223301CB4CB4984800000004DA40101A0990D90860C1830494";
    attribute INIT_3C of inst : label is "14545155115115115514545151155199991111999117DF7DDFDDDF77DDF77F7D";
    attribute INIT_3D of inst : label is "02030020F8020212ACE85C0E84AB3A570384B2C84B6C9BFABEEF675475D15515";
    attribute INIT_3E of inst : label is "00210040040000002041040100081090000502428000000440D0824480030080";
    attribute INIT_3F of inst : label is "38D041100912102408034410482202800020082942121008282C3401A6000C20";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "005838034014AD5AB56A4489122D5AB56A4489122D5AB56A960D1896AC4876C1";
    attribute INIT_01 of inst : label is "2EC0BC57AAED485932716AB402C248E892490482492490A4D48A91526A4D4897";
    attribute INIT_02 of inst : label is "0410101CEBB0028AD7EBB5063CC724AAB2324664CC7012D0824001884084222F";
    attribute INIT_03 of inst : label is "9C14C99A487253921C90E4A7243921C9464A3241928C9460A3288CA080830001";
    attribute INIT_04 of inst : label is "9D59AC5C1449C1449C1441C1441D172A4A02A0A0C14C9C14C9C14C1C14C1C14C";
    attribute INIT_05 of inst : label is "888A9586A5596435645965116511403E8E208374099AE942ACA49224591A774A";
    attribute INIT_06 of inst : label is "05A51160609281D6D11688B2884D49A64A46594459444A2157229AAA22A71513";
    attribute INIT_07 of inst : label is "0E14F0A3A51C29E9468ACC6E1508242455CC020B0414400C80110430494092C1";
    attribute INIT_08 of inst : label is "3829B043160A6260E3261D29E94F0A3AD18816601660E7071831C1864C307393";
    attribute INIT_09 of inst : label is "66495EC3429508160208158C92DB04100459294E729E086C10C58218F0531324";
    attribute INIT_0A of inst : label is "0404095011244492A99355931F063831C9C55449448892553262C18D4A4E6354";
    attribute INIT_0B of inst : label is "84142C8A4E60B35C0A084C8B3073D4E2124A869322CC18F5704201950D5042DD";
    attribute INIT_0C of inst : label is "00EA982F1249219939E0424354B660C78482168C0214AB25912D921400CB2E88";
    attribute INIT_0D of inst : label is "06966596DEDB5511CB459B1D0DDAC624B9768B2D500B04C61881D99999D8154B";
    attribute INIT_0E of inst : label is "8EAA60B4D47516161564A39B720A9D700D965B6A9A61166C0308B2C36D16DAA1";
    attribute INIT_0F of inst : label is "C731E4D556ACA032EC8CBB84277D30B00ADA85A4A411B486A16C52900105CEBC";
    attribute INIT_10 of inst : label is "A8EC9E10471C71C71C70C30A25D7115061C78E625D092CF03C225B9CD7399CEE";
    attribute INIT_11 of inst : label is "A33400688AC0D048340520C0803E8E2158DCBCF0E2E735CE6733CB1CC7393555";
    attribute INIT_12 of inst : label is "B4B241830C1C64C3271830C9C78C0020B60D15F4C7AE3D30E986B061EB4A0E30";
    attribute INIT_13 of inst : label is "BE5F9CD9126B2DC42E0A2C632ED8FB05B83961C71C71C71C71C71ABA83506341";
    attribute INIT_14 of inst : label is "239D1091AA892B510B5101019248A351CBAB1D52A34BEAA34DBEDAAA4BEAA34D";
    attribute INIT_15 of inst : label is "3044C214F517AA4C8040ECC0C9D98322E8DD91C4E84922C6C9319BE441F42492";
    attribute INIT_16 of inst : label is "6D5ED8982B5ED94C11AF6CA608D7B653046BDB2982B5ED94C15AF6CA60AD7B65";
    attribute INIT_17 of inst : label is "B2B2D8CA927C6D564E19B31D8C6CC531B1D9A7677FF7F46929270A71B754DBAA";
    attribute INIT_18 of inst : label is "000000001008286D8204004083430A000090C00000084004B1D95436C6DEF272";
    attribute INIT_19 of inst : label is "1041001041001041001001040000092A60004284C010080002CA0A94040000A6";
    attribute INIT_1A of inst : label is "0410410400410400410400410400400410410100104100104100100104104100";
    attribute INIT_1B of inst : label is "8DCAFEA0002B735314E6AA7151068105B7140036D17CAA040041040041041041";
    attribute INIT_1C of inst : label is "B3BA048005912856E520A18005E9525027794918A04586CA1453008885155491";
    attribute INIT_1D of inst : label is "2567283840B25B08252C049465564958A22D0645F2A35120B951A84A9504E6AA";
    attribute INIT_1E of inst : label is "0000000000000000000000F420B4E04C9A023987090D4B48840009400502C250";
    attribute INIT_1F of inst : label is "000001FFFFFFFFFFFF21043FF800000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "08100081000804008033FFFFF8CB008E029405382A5C01FFE001C01FFFFFFFFE";
    attribute INIT_21 of inst : label is "0004404242040446068040080810008100081000810008100081000810008100";
    attribute INIT_22 of inst : label is "4E64125790911991111088088880155555821A6846901141800007FFFFE00000";
    attribute INIT_23 of inst : label is "0CB4A624402839030912DEC64941E83C80446804124004124100811CA1669583";
    attribute INIT_24 of inst : label is "B2B25860B2B2C3463A40021200021A40021200020804B64B64A4B64B64AD28C3";
    attribute INIT_25 of inst : label is "9649AD2974A7A51C28E1461A2CACB0C16CAC961830D1868C3461A30D1868C305";
    attribute INIT_26 of inst : label is "0085394AD694E5CA800087294AD694E5DA400087394AD694E5CA002828281600";
    attribute INIT_27 of inst : label is "D694E5DA000085394AD694E5CAC00085394AD694E5CA800087294AD694E5DAC0";
    attribute INIT_28 of inst : label is "82008539CAD694E5CA42008539CAD694E5DA00008539CAD694E5CA400085394A";
    attribute INIT_29 of inst : label is "87843C60E307083841C21E10F1838C108539CAD694E5DAC2008539CAD694E5CA";
    attribute INIT_2A of inst : label is "12D9D21E90F487843C21E10F487A41C20E107083A41D20E9071838C1C20E1070";
    attribute INIT_2B of inst : label is "0080000000040000804703880430308040000804000081C0FC0E3C0FC0F1B5DB";
    attribute INIT_2C of inst : label is "61895ACA0100FA3881BC0FC0F1C0FC0E04000080400008043030804703880400";
    attribute INIT_2D of inst : label is "0562C2D46AC02F10C4009842C06AC158B0B51AB00BC43100D6280100C00496C8";
    attribute INIT_2E of inst : label is "2A9ADCEF38822C415822208A6B33BCE208B104608A35D7B06D2CACCEB855A8CB";
    attribute INIT_2F of inst : label is "882B339C6208B104608A8A21ADCE718922C41582AA2AA6B73BCE248B10560A88";
    attribute INIT_30 of inst : label is "848885BB801B8EED00371DC512B6801B8ADC00DC771112CB34E25491A470F4A0";
    attribute INIT_31 of inst : label is "C43E01F007C05F017C04B64C6F5E3C561C9880D248A0B425505A12A80D091406";
    attribute INIT_32 of inst : label is "0EA080498C96C44A4CA1C2A900BC9596B6D6CAC954E60315AD69A2F8F7CC2424";
    attribute INIT_33 of inst : label is "D7CE1AB800568294C3096CA40100C13044109FB406798C4949073C025B2B742D";
    attribute INIT_34 of inst : label is "64C26AE64697CC98DD880C4127349A40004071F8E3D036F332D8EBCE40870028";
    attribute INIT_35 of inst : label is "E4C6D5D3FFE0007333300C2D2CE60B34B8B32EDA6599923149999D99CF23CB39";
    attribute INIT_36 of inst : label is "4C91003B801BA76801BA744596D00374B7003748EE8CB36DCB9693D0C6C86E0E";
    attribute INIT_37 of inst : label is "BC4B12048191838306432648A1932450C992A864C95432648A1932550C992286";
    attribute INIT_38 of inst : label is "D2FD987338C18C2D25E82B659603116A3124DC580CB51A66399C60C616D2FD9A";
    attribute INIT_39 of inst : label is "0814C20015A87338C1882DA5E82B65960311603124DC580CB01A66399C60C416";
    attribute INIT_3A of inst : label is "BDB5B5AC96C9ADA2800AAAA0002AA802800492EF01C4DC9B88425380AF639813";
    attribute INIT_3B of inst : label is "5755E333323333323250D555550D31CC804C9B7300063D03B8EA18E3468D19BD";
    attribute INIT_3C of inst : label is "450514015415415401450514144111911199119919355D5F55F757D5F57D5D5F";
    attribute INIT_3D of inst : label is "E54CDA01F47102128CC1C83C84A330320F04A4104A010625E9198CDECC641141";
    attribute INIT_3E of inst : label is "52F4EB0B1AB53D65D1A242CCF33E5C7D7BA187E148B1EF9EB4DD61B767A5E333";
    attribute INIT_3F of inst : label is "11555E55471E2E3C59E3DC5C70E107185800D0BB885ABAA0D191B370D3CD53A4";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "556602AA316F9FBF5AB5FBF5AB5FBF5AB5FBF5AB5FBF5AB457F81AFD2D788C0A";
    attribute INIT_01 of inst : label is "BBDF2AE7C3BE2A7DEAD5EF33BC8EC0F9F5BAFD6CBE5B2F5F6BFD7D8FF1F63FD0";
    attribute INIT_02 of inst : label is "8EEAC8E70302A4FA8621F44707B610113E9B3736694BBE2B8948CD63717038A9";
    attribute INIT_03 of inst : label is "F91437F48A444222111408A044032011088A44522211948C808806F75662EEAC";
    attribute INIT_04 of inst : label is "184D0E7914BF914B7914BF914B715F8C2318C230914BF914B7914BF914379143";
    attribute INIT_05 of inst : label is "2A038329110011481100114811001B8C5551DE47DD5CB84120138A142B74E581";
    attribute INIT_06 of inst : label is "4D914814A4D542C11008800880A32A20854206400440220187E1EFF38A3A57D9";
    attribute INIT_07 of inst : label is "931418A0ED27213108027B4370BA36B7C180249B6D36934D269369A49A49349B";
    attribute INIT_08 of inst : label is "2321664294C8534DE44607213909980E406CF35CF348C046033819C0DE467223";
    attribute INIT_09 of inst : label is "33670D948E76FB731E7AF03A6D36B6C93DADCE77B08C8A5910A52214A4529E64";
    attribute INIT_0A of inst : label is "1B6387084EDDD0582D5A25338267023811CA63AD3BBA0B05AB4C99C26F6B5A1A";
    attribute INIT_0B of inst : label is "7CF3E6B88E138A14948077F9A66027FC7465201DFE69980875DE240A00200322";
    attribute INIT_0C of inst : label is "58FFCC2F1DC738D23819C3F4139B4CE067DE9BB59EF797BCCCE6DDF16C6A3C3B";
    attribute INIT_0D of inst : label is "9BDB34D24A49E516ADF1C3BB0F1D80C0D1A7E38EEAB258CD38EC9C9C9C9FBAB2";
    attribute INIT_0E of inst : label is "29FF30BBFF5FD85856C3E1C92DDFDA45CCD3493C9E76470EE3B238E127124F21";
    attribute INIT_0F of inst : label is "5CF5ABDFE4B549DF3677CD7CE9A6752F1554FDC450018A001F29461CF76F242A";
    attribute INIT_10 of inst : label is "32B6835C9451441041051454492C7246707293DA950794C8B23FCE7EFCFDF3CB";
    attribute INIT_11 of inst : label is "9BE8017F4C6FA4B4699CD1B79B8C5550DEE3629DE79FB73D7CFA6D73D5AEF7F9";
    attribute INIT_12 of inst : label is "69264223119C88E446023811C26A604AA102011CA0E507293B40266043F8CC17";
    attribute INIT_13 of inst : label is "E97ED6AD7519E690BD1889E93BC68247F4F69F945145145104104425504670CB";
    attribute INIT_14 of inst : label is "5AF5AAADFF2DB09010901E2224930A878240F00B9AEE839AEBE9FAC1EE838AEB";
    attribute INIT_15 of inst : label is "60E7978781471FD852C314EEA629BA95A5344A5243DD959FA4E7CEB577A1EEC9";
    attribute INIT_16 of inst : label is "2E9B57307A9B5698394D8B4C1EA6C5A60F5362D30721B16983D0D8B4C1E86C5A";
    attribute INIT_17 of inst : label is "949568527BE4B4A97A0C99DC8464651190C8A325E8208158532D5CDCB3FE59FF";
    attribute INIT_18 of inst : label is "00041001017653E2128009F49F1CD4E0223DE8800000041FD0CA25125B4C6A02";
    attribute INIT_19 of inst : label is "124124124120124120120120DE3E364FD108070E27D108137DC5D3F7DD80837B";
    attribute INIT_1A of inst : label is "0480480480490490490480490480480480485120124120124120120120120120";
    attribute INIT_1B of inst : label is "28EDDD4F5502287A8D50832A7A9B9C50E2A78A1B72F48B848049048048048048";
    attribute INIT_1C of inst : label is "E4D02EBE0B22EEBF77C1BABE0BF32291F5FA157202EBB8D3AB9E1AD5EAC1E157";
    attribute INIT_1D of inst : label is "D410A3021909444314C0E050940885006A59444BAA1D0F28D50E8753F5DF5483";
    attribute INIT_1E of inst : label is "020040000042000004000361CA8115234044061CA4421C1132B4251848241140";
    attribute INIT_1F of inst : label is "0000000000000000004040B807C000020020024000006A002104000200210400";
    attribute INIT_20 of inst : label is "600006000066638D74C80000030100707050E0A1C14000300000000300000000";
    attribute INIT_21 of inst : label is "0000000000000000002638D70008060080600806008060080600806008060080";
    attribute INIT_22 of inst : label is "B9FA9F98E2BF77777FFFEE666EC015540014041010520C104007F807E01FE030";
    attribute INIT_23 of inst : label is "49A2299116454CADB4C9B7BF24AB654DB495B241949A6D2650453635CBA32E9B";
    attribute INIT_24 of inst : label is "0584B27821A19381A204041414140205051414140E5A69A69A3A69A69A31CC92";
    attribute INIT_25 of inst : label is "C9A529085CE4E7063831809E086864E001612C9E04E027013809C04E02781380";
    attribute INIT_26 of inst : label is "4A99DEE798E7796C184A99DEE798E7796C184A99DEE398E7796C1877622264AA";
    attribute INIT_27 of inst : label is "B9E7796C184A99DEE7B9E7796C184A99DEE7B8E7797C184A99DEE7B8E7797C18";
    attribute INIT_28 of inst : label is "184A99DE67B9EF797C184B99DE67B9EF797C1A4B99DE67B9EF796C1A4A99DEE7";
    attribute INIT_29 of inst : label is "E0C7067833C19E0C7263833C19E0CF0A99DE67B9EF796C184A99DE67B9EF796C";
    attribute INIT_2A of inst : label is "C9B773931C9CE0C7073831C18E0C7263939C98E4E7263839C19E0CF067831C98";
    attribute INIT_2B of inst : label is "6D5EADB6DDEADB6D5EA8B455EA8B455EADB6D5EADB6D5C2D02D0C2D02D0D2D55";
    attribute INIT_2C of inst : label is "D3B4F333186E31554642D02D0C2D02D0EADB6D5EADB6D5EA8B455EA8B455EADB";
    attribute INIT_2D of inst : label is "2CEAE73836D4F175E16D26672836CB7AB9CF0DB51C5D785B17B3609D6E674D31";
    attribute INIT_2E of inst : label is "B324E0B8F332E333933A0CEC93C2E3CC8B8CCF4CCA177952BA3F4F0B067E707B";
    attribute INIT_2F of inst : label is "EC9382C34C8B8ECE4ECA3B334F0B0D332E3B3D33A0CEED3C2E3CC8B8ECF4CCA3";
    attribute INIT_30 of inst : label is "FDCB879135A9BE446B537CDFDF9A35A9BA69AD4DF375DE79ED86E7BD6E43C38C";
    attribute INIT_31 of inst : label is "58C9984C6131C4C61319B6C66C58D1A979F1643CDCD98FEF6C87F73663FBDB21";
    attribute INIT_32 of inst : label is "4C7B7DAEAE4D9DE5668D8CA7CB0FC3DC7F0F71FE17ABBDB735CF419ACDCFBFEC";
    attribute INIT_33 of inst : label is "6C547C92B557FE4534F4D33964599745996762C9FB9237FECF7DF1CD34CC5FE2";
    attribute INIT_34 of inst : label is "69973EECEFF3D98CD4DB06C063363EC07F890E90F9A93EE43AEAF12FA57E5AAD";
    attribute INIT_35 of inst : label is "6C66E5B7555555311119C28B36722B19B2BB35DA65C9F31B9888898CE651BB19";
    attribute INIT_36 of inst : label is "C7B9B9913599B223599B3675F346B3349A6B3353E6EAB9A5DCDB72DBCAF659D3";
    attribute INIT_37 of inst : label is "BC771FDDA5A5B7A7B9B363DED9B1EE6CD8F7B66C7B9B363DED9B1EE6CD8F7B66";
    attribute INIT_38 of inst : label is "F2FD999750B9FDEBE5AEE6E5F9E17794176C4FE787CA0EE5A3E85CFEF5B2ED9C";
    attribute INIT_39 of inst : label is "1FA4D8AD55FD9F50B9F9EB65AEE6E5F9C1779C176C4FE707CE0EE5A3E85CFCF5";
    attribute INIT_3A of inst : label is "474E4E334D36782280A0AA0A0A8002A83CB7E98A5BCBF58999CE332BDF479DF6";
    attribute INIT_3B of inst : label is "81D8B3B2233BB2233B28E1E61E0AA17744661235291B58E4D6C4A16FDFB76F67";
    attribute INIT_3C of inst : label is "0EC45143BB11B11143AEC45B10B1599D91911191599D8BD88189F6209F620BD8";
    attribute INIT_3D of inst : label is "38A022DC62AA8FC99EAA656DF267AAD95372E9372ED27368BA4D355554CB15B1";
    attribute INIT_3E of inst : label is "00A0C000AC4880AA29D024AC2078902143C210C00781C679325303061E511941";
    attribute INIT_3F of inst : label is "174C288628910142864E2A331CFB51DE8E0F0306B0930343260241A1612C944A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "D43426A1A067B264C993264C993B76EDDBB76EDDBB76EDDA3EB986ECC373DCC1";
    attribute INIT_01 of inst : label is "D9938372E1930471E1C1C7869E5EC8F9B1D8EC7633198CF7FEFFDFFBBF77EEDC";
    attribute INIT_02 of inst : label is "C6798C13A1301E6FC3ACB440621A06838ECD839B33199E678739CCF7B3781CD1";
    attribute INIT_03 of inst : label is "E1018E2080C41620B105880C406202101882C41620B101080CCA4233CC666798";
    attribute INIT_04 of inst : label is "166C8461018E1018E1018E1018E0198C6318C6301018E1018E1018E1018E1018";
    attribute INIT_05 of inst : label is "6339932D906D906D906D91499949BBE0FFBFB5FD83BEA985A7D24D9325A4754C";
    attribute INIT_06 of inst : label is "6C116D9100E84419048824CC247B230DB118641B641B30D8C3E3E557987AD2BD";
    attribute INIT_07 of inst : label is "2101080C40420210100121B17439B9BBD08624906DB2DB6134C249149A0DB65B";
    attribute INIT_08 of inst : label is "420A0414108283880C406203101880840633F30BF3080840620B105080840420";
    attribute INIT_09 of inst : label is "398F4996DE72B9F12C78F67B69361249BD0C84A12C6080C10184203084061C40";
    attribute INIT_0A of inst : label is "1B0A4F664ED9D8EC8E1C7820A040620A10105B6E3B7B1D99C3AF101A71710D9E";
    attribute INIT_0B of inst : label is "3C59E67882879D019624B3398416678EF325892CDE61059C03DE67631B31B5B3";
    attribute INIT_0C of inst : label is "D0D55B2D1E6592C2033BC39E5F8B0808E71E1C319EF3343C49E2C6F33E613B79";
    attribute INIT_0D of inst : label is "5CDD71C6D8DB76370E31C3720E1D8368E1C6638D013AD4F928E59D9D9D9C003A";
    attribute INIT_0E of inst : label is "03556CB9AB2ACCCCCB83425B68005F6D0DC71B6EDC6CC70D936638DB6E06DBB3";
    attribute INIT_0F of inst : label is "4DEB27AABE1B69CD9A73663DECD6C5BD0FB6BC63186C630D8F04129D7F6FE60E";
    attribute INIT_10 of inst : label is "96371340BCF3CF3CF3CF3CF6482456440620210CD600C05E1793D6F4EDE9F3A4";
    attribute INIT_11 of inst : label is "8CC86161417120B44CFCD137BBE0FFBFC2E7464005BD3B7A7CE96137AD89EAAF";
    attribute INIT_12 of inst : label is "420404203105882841420A101A64035ABD030EC80C406203101A0416207882C7";
    attribute INIT_13 of inst : label is "C364C66C73D9C7B03111FB81B1364EC0C7C3BE38E38E38E38E38E60446440692";
    attribute INIT_14 of inst : label is "CC4AC74155F5DCD6DCD6DB1B2492856E324CC7511D84391980C3652A84391980";
    attribute INIT_15 of inst : label is "66F7337B1EB2DFD813871CCE6639B99F27E4DAD6B7D6CD9D366F6C1B8F5BEB6C";
    attribute INIT_16 of inst : label is "6F9BD3B37B9BD259BDCDE92CDEE6F4966E737A4B3739BD259BDCDE92CDEE6F49";
    attribute INIT_17 of inst : label is "CECCD83A06D36C56D90DB10E4CF2CD33C9E5A7980A80AB94D36DDEDDB6AADB55";
    attribute INIT_18 of inst : label is "0000000000473232820000DAED90EC8000B660040000408D89E63716F6D8C81F";
    attribute INIT_19 of inst : label is "10410010410410410410410068802C682008401174100001A46B1A0042000108";
    attribute INIT_1A of inst : label is "0400400410410400410410410410410400400104104104104104104100100104";
    attribute INIT_1B of inst : label is "02206A8904098A18D314008818C36514C880A29B6CB501041040040040040040";
    attribute INIT_1C of inst : label is "080BB108004002031000080800C002D05A8F6240BB10CA6081D1166E20441624";
    attribute INIT_1D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFBFFFE88AB2D3564CAE565A66572B5A01411408";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFE000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "F7EFFF7EFFFFFFFFFFFE000007FFFFFDFDFBFBF7F7E3FE001FFE3FE000000001";
    attribute INIT_21 of inst : label is "000000020240004202FFFFFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFFF7EFF";
    attribute INIT_22 of inst : label is "D198DD8C70AE6EEEEEEEEE6EEEF02AAAA977D77CF1C75C77C3FFFFFFFFFFFFC0";
    attribute INIT_23 of inst : label is "450209110764408C366D2119B62A256536D78024804800920924172460D18343";
    attribute INIT_24 of inst : label is "4849020B6C6C1010D20200100200120301100200161B4924925B492492588410";
    attribute INIT_25 of inst : label is "6DB25A96880C406202101882D2120416DB1B6080841620A105082C416202101A";
    attribute INIT_26 of inst : label is "1258D63108431826181258D63108431826581258D63108431826180888A275A3";
    attribute INIT_27 of inst : label is "08431826181258C63108431826581258C63108431826181258D6310843182658";
    attribute INIT_28 of inst : label is "181218C63108431826581258C63108431826181258C63108431826581258C631";
    attribute INIT_29 of inst : label is "6C43621B10D086843421A10D086C436218C63108431826581218C63108431826";
    attribute INIT_2A of inst : label is "ED2621B10D886C43621A10D886C43621B10D086C43621B10D886843421B10D88";
    attribute INIT_2B of inst : label is "92215249221124922110482211448A2112492211249222120121012012066274";
    attribute INIT_2C of inst : label is "21B6A1207DEF83FEF8012012021201211124922112492211448A211048221124";
    attribute INIT_2D of inst : label is "A1C2CB602CF0F81B236266CB602CE870B2D80B3C3E06C8D857BB607DBCDF6923";
    attribute INIT_2E of inst : label is "3322E1D8E7A0C78B93B29CCC8B87639E831E2E4ECA130D50D83B2F1C66C6C063";
    attribute INIT_2F of inst : label is "EECBC7639EC31E2F4EEA73BA2E1D8E7A0C78B93B29CCC8B87639E831E2E4ECA7";
    attribute INIT_30 of inst : label is "25CF87367173F0D8E2E7E1F81C367173F0DB8B9F87E11CE3DDB2E4B92E5F1F1E";
    attribute INIT_31 of inst : label is "79D97CC8F3238C8E323930C42C5B870BE0C66425DC99092E4C849726424B9321";
    attribute INIT_32 of inst : label is "EC4079860F691BB1B35E4C2EC30B6168290520A6474398A97A5E4084C42F9F8C";
    attribute INIT_33 of inst : label is "D98A0EB6AC173E4126769258F63D0E4390E3305BF9D6B2760E3CE7EDA4960FE6";
    attribute INIT_34 of inst : label is "65D774CCCF23198868F347836218B2C00000000013A83A2D3EF473C66338D60C";
    attribute INIT_35 of inst : label is "8C42C59600000161111F9A3E7AD69B10B2BE78DFC5D8671BD888898DAED30B11";
    attribute INIT_36 of inst : label is "C4B9FBB6715BF6C715BF7D0586CE2B7E36E2B7FB0F88B3CDDE5CEB473CE659D9";
    attribute INIT_37 of inst : label is "B4791C5966666464DC32625E99312F4C9897264C4B932625C99312E4C9897264";
    attribute INIT_38 of inst : label is "66C9B64D2863C3C64DDFCA0DDB01E5B01E6E5D6C06D8082E109431E1E366C9B6";
    attribute INIT_39 of inst : label is "0534F1AB05C2452863C3C6CDDFCA0DDB01E5B01E6E5D6C06D8082E109431E1E3";
    attribute INIT_3A of inst : label is "6363631B692318B5FF55F5FF5F5F5F5F5C33F5AADD2F6188C4210B6B05C099E6";
    attribute INIT_3B of inst : label is "7DF7D000000000001150141141050000000000638009E4766646339FBF7EFF63";
    attribute INIT_3C of inst : label is "4141454045045045404141450450408888888800001F7DFD7FD57F5FD7F5FDFD";
    attribute INIT_3D of inst : label is "71F0E1DF07FDFDEC0B2205457B02C8C1597B49A7B4DB754D5355567567450450";
    attribute INIT_3E of inst : label is "FEBC3F8FF7E7E7A6BD7A7EF5D7AF4FCF3D38FD78FF1F79E3AF5C7D3A71F8FD7C";
    attribute INIT_3F of inst : label is "D34F35D335EBEBD3CF9D63F1CF3CFA63F79FD3A6B8EBEBF9D3D3D63E9A7BF7E4";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "7C1223E010228912244891224480000000000000000000007E3802AC01534C03";
    attribute INIT_01 of inst : label is "48B90720C0862450A9414503940A48C89148A45229148A16A2D45A8B516A2D4C";
    attribute INIT_02 of inst : label is "863888568100B42F82A534C1263200111A44A28913188A628F7BC6C631691541";
    attribute INIT_03 of inst : label is "43048401824C026013009804C026093009824C126093049821880631C4426388";
    attribute INIT_04 of inst : label is "126C044304843048430484304846118C6318C630304843048430484304843048";
    attribute INIT_05 of inst : label is "212497003000B024B000B100B1008000000137998A2640C72753499325A47215";
    attribute INIT_06 of inst : label is "003100B010A1C04B001800580069610497092C092C09604983A125548A4852A4";
    attribute INIT_07 of inst : label is "83041820C126093040036313D0E9A9AB40800001249049209241249241200000";
    attribute INIT_08 of inst : label is "26000C001180029820C126083041824C1063530B531820C106003009824C1260";
    attribute INIT_09 of inst : label is "20050B801AD7EBD37C2852692480B6DB14AC421080018203040460808C1014C1";
    attribute INIT_0A of inst : label is "094E45224A4B48A48A14226094C1060830405B6A29691491428430405353189E";
    attribute INIT_0B of inst : label is "14CCA66182129C019C0011698C1062A6536700045A630418015A6D2E09609096";
    attribute INIT_0C of inst : label is "50554A651A2CB6C60139429A4E9B1804C50A15398AD73C14D8A6CE537A61296B";
    attribute INIT_0D of inst : label is "505128A2484946940868A972060F83088102D1440430506828D4CCCCCCCC0030";
    attribute INIT_0E of inst : label is "0355299B2A8AA0A0AA8342492AAACE2544A28928CD2DA2A5B96D145926024A39";
    attribute INIT_0F of inst : label is "04A2028ABA4929448A512215845245B50E92152170242E0485010424354A2202";
    attribute INIT_10 of inst : label is "923211C0B0C30C30C30C30C2586CD24C00608318C85450C8323152D4A5A956A4";
    attribute INIT_11 of inst : label is "99806141213000BC05D4F01680000000C2A3424044B5296A55A920128880A2AE";
    attribute INIT_12 of inst : label is "090C026083001804C02601300A200A0A1F060CD820C1060830400C1000298202";
    attribute INIT_13 of inst : label is "8144436CD34983142300F108A0320C408282B434D34D34D34D34D20DC24C0008";
    attribute INIT_14 of inst : label is "58C8850155D55580158019022493852416444200080010080081440000100800";
    attribute INIT_15 of inst : label is "64C63142382257580B873C995679655D07A0D6B5955A54B512AD2428854AAD25";
    attribute INIT_16 of inst : label is "260B13326A0B12193505890C9A82C4864D41624326A0B12193105890C9882C48";
    attribute INIT_17 of inst : label is "CC4C483012532406490C911A4652641948A482980AAA010442259EDC92AA4955";
    attribute INIT_18 of inst : label is "00000000102C323602004002AD918C80008020002100000008A623127248581F";
    attribute INIT_19 of inst : label is "10410010410410410410410420120D42000040816010000092EB50914000108C";
    attribute INIT_1A of inst : label is "0410410410410400410410410410410410410104104104104104104104104104";
    attribute INIT_1B of inst : label is "032228294509CA1A139409C81A036514DC80821B649408041041041041041041";
    attribute INIT_1C of inst : label is "9A21150804D126139120980804E8108058062A50115448298580060E614042A5";
    attribute INIT_1D of inst : label is "000000000000000000000000000000089BB6C156D6AF56D82B57AB1090439000";
    attribute INIT_1E of inst : label is "FE007E42427E007E060202000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "00000000000000000000003FFFE10A52A528427E4A4A6E003FA723FE003FA723";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0102500440AEE6666666EEE66EC8155554800001040800800000000000000000";
    attribute INIT_23 of inst : label is "00160030950C05849080003000E10C0012160124100020824924040001400502";
    attribute INIT_24 of inst : label is "0000060124243009910200100200110301110200000000000000000000001000";
    attribute INIT_25 of inst : label is "008542509820C1060930418000000C02490921804C106083041824C126093040";
    attribute INIT_26 of inst : label is "3200121084210860003200121084210860003200121084210860000A0A2860A0";
    attribute INIT_27 of inst : label is "8421086000320012108421086000320012108421086000320012108421086000";
    attribute INIT_28 of inst : label is "0032001210842108600032001210842108600032001210842108600032001210";
    attribute INIT_29 of inst : label is "24C126083049820C106083041824C10200121084210860003200121084210860";
    attribute INIT_2A of inst : label is "80026083049820C106093049824C126083049824C106093041824C1060930498";
    attribute INIT_2B of inst : label is "0000000000000000000000000040080000000000000002000001000000042015";
    attribute INIT_2C of inst : label is "9112949050000000000000000200000100000000000000004008000000000000";
    attribute INIT_2D of inst : label is "00C24B60264048120142664B6026403092D8099012048050F2A900513AD52492";
    attribute INIT_2E of inst : label is "A20244C086918603162A1A880913021A46180C58A81004C04220244C6646C049";
    attribute INIT_2F of inst : label is "880913021A46180C58A86A20244C086918603162A1A880913021A46180C58A86";
    attribute INIT_30 of inst : label is "218E041A2151C06842A380E014142151C0510A8E038114415DB0C4310C5A0A1A";
    attribute INIT_31 of inst : label is "75D950C843210C84321112C4644B063B408250649894190C4A0C862506431283";
    attribute INIT_32 of inst : label is "EC8260A208002885C00800280109212424849090440401A98A6240C84646022C";
    attribute INIT_33 of inst : label is "998A1422A8323AC002D2490842108421084550DBE14290508815A3A492421FA6";
    attribute INIT_34 of inst : label is "21873E6ECC235D88C8E1470B623030C000000000196018441A54D1CC21105418";
    attribute INIT_35 of inst : label is "2C46448600000121111F5E3E2A528918969F28CFC4C8831BD888888CA4510911";
    attribute INIT_36 of inst : label is "C431EB9A2149D342149D39048284293A144293B007089104D8500A022C655900";
    attribute INIT_37 of inst : label is "946918F160606060512B621895B10C4AD886256C4312B621895B10C4AD886256";
    attribute INIT_38 of inst : label is "325C924628410686E4C38B24DB01C5B01C6C496C06D808461114208343325C97";
    attribute INIT_39 of inst : label is "082040AA0C82462841068664C38B24DB01C5B01C6C496C06D808461114208343";
    attribute INIT_3A of inst : label is "000000092494180A0228888222088A20B0004188540A25884842112A20C209C6";
    attribute INIT_3B of inst : label is "FD5FC0000000000011616666661600000000007C000B00F00240020891224400";
    attribute INIT_3C of inst : label is "40155510005405551000154054054088888888888895FD57FD7D55FFD55FFD57";
    attribute INIT_3D of inst : label is "9815360000000D8008602C216002184B00600096004875715C5541F41F405405";
    attribute INIT_3E of inst : label is "038500C070A0A0A2850A0A9554A951534B4D050A81A74C34A946050A980C070A";
    attribute INIT_3F of inst : label is "554714531C3A387468C5703AE9868A3054C050ABAD38382A70705282AA3A7466";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
