-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "D352A0B17FEA2A4977BB18080082410493A07FF3F4CB65F5D87EA7A3D3F3EAB0";
    attribute INIT_01 of inst : label is "208B53050688596AA28094500A24F28449614EA8FBC4F2612971B05C07AC02D0";
    attribute INIT_02 of inst : label is "FC616582249E4F061E45A982F79FCB31445F3FC419F84F3FD72089804BBC4109";
    attribute INIT_03 of inst : label is "89BE341034499CAFCD9900410F7AFFA7DC55555E004169FD4262E38A88145499";
    attribute INIT_04 of inst : label is "51A089270943A937ABA93780076A8522A21166842AD64C1728AB834409386F50";
    attribute INIT_05 of inst : label is "F34F2110D2108910805499B883E2D415122286315425C47E8BC50155075D544E";
    attribute INIT_06 of inst : label is "4250545C51EB4B32A602B64FB4BA4DFDB349E496C9BD51493C0A4D0060F24174";
    attribute INIT_07 of inst : label is "829D5134F22CF4224501505499A48FD17E8F9C5A14936A1964B0AAA294A2545C";
    attribute INIT_08 of inst : label is "830615560605408A9137523A1328A7118145084A0E87140824D26D52CB94E216";
    attribute INIT_09 of inst : label is "54CA121CA721674943381D902702F8AD58C58A4236918946074DE28A00013802";
    attribute INIT_0A of inst : label is "0124C9D65DF6D4EBED1FB80AFE698E58E7331252C1201AA28426A43896244542";
    attribute INIT_0B of inst : label is "E5EB397467B396ACE5D199110A51D6846A3DD99A0867819214870E9F122A1D48";
    attribute INIT_0C of inst : label is "6B64AA0978053234FBB84E2BE5E79653807D913E85137D246FA142D79E5651EC";
    attribute INIT_0D of inst : label is "0065F669E00041882DCCBD13E898CBF13E89886EA5A11A3AD6B1955958B5A7F2";
    attribute INIT_0E of inst : label is "85B548468F01009124598E6A22882AD59ADD56D23D4A4ED952BA0284EDB65400";
    attribute INIT_0F of inst : label is "F4A295C73B654AE89C589DB05B731885559263340305B27CBA5FD229C587F434";
    attribute INIT_10 of inst : label is "27D74148A8F2CCD0C9353354A479EDB68DB55592F44F98D5564BF13E621BA97F";
    attribute INIT_11 of inst : label is "EF7F119E3768C5EE6CFBDFF11A5D76E27AF816A69B46E37D78F97539621AC572";
    attribute INIT_12 of inst : label is "0B1A0B4450962510C48201547BBC4D10C674809C06DA3A2A108350F7389A30C4";
    attribute INIT_13 of inst : label is "484546A0EB0C9838679E65AF8E3E72652C5C8E34B5E45FD06081452A445AAA44";
    attribute INIT_14 of inst : label is "8D091895221247ACE12504A77646438F3932923D66776324EA4B7A2164EB4C15";
    attribute INIT_15 of inst : label is "8BC8E48A2FFFFEAA720B26212262E221589B4358CA17429C88993C46D35C0290";
    attribute INIT_16 of inst : label is "B3CF40838708A302315814F5635D52D15505BA343741AA2A41A13CB261A14808";
    attribute INIT_17 of inst : label is "A88551C7AA801570B00337378DF741A66D0AF7DBC646754A7661364651397DDF";
    attribute INIT_18 of inst : label is "06845ADA168B448DC8AA48A4CCE8D70C5F2D812B88F7399A39CD38191D296092";
    attribute INIT_19 of inst : label is "2E7BFF822726DCCCE49B8C34294A3110D7DC0BC7E82692858267E886AC18A310";
    attribute INIT_1A of inst : label is "51100284406842221250C068413219260C34CC01030D25967F30100000C02B02";
    attribute INIT_1B of inst : label is "23203282323242020440010427986DFAC27C11028CBAFEA0114670009ED2FE3D";
    attribute INIT_1C of inst : label is "0A78EF5A24BC64930D0D10402032C320EC4A2C458A8D5406EC19E94100801669";
    attribute INIT_1D of inst : label is "00000009C4060000F640080036401F003654204404AD120482E8110842108421";
    attribute INIT_1E of inst : label is "4A5569652AAAACD345656565655559EA9EAD555575DD9E6EEBAAAEBB9B6775D5";
    attribute INIT_1F of inst : label is "037C32C8EAFDF2A94008E2C01A112E6B985A1681AA680632A8755570AA74D6A1";
    attribute INIT_20 of inst : label is "7BF7A77B4826D648F836A54A89FFC719E08ED558FD7FC8763CABA0288D3AA281";
    attribute INIT_21 of inst : label is "994F3A2F708DAA1734B67BEF3EE807D75DF787E687CB6FC2577BEBD43C25B01E";
    attribute INIT_22 of inst : label is "75537C2090000154D0D151EA3B56A3D92E0B48F8B7CFC9E23418CA7F49226965";
    attribute INIT_23 of inst : label is "EF6A66D01B99AA2BEE638E1870A4299A9E2222FDDD71749C679F44EAA312E843";
    attribute INIT_24 of inst : label is "C40C0048CF0481103A36F19EA8A0800D0404680003400118234E7B5997FE934A";
    attribute INIT_25 of inst : label is "2224F385852C020192E181E4CDA07F3FDCF4FE196E9E0F6E87C0E8012A3517C6";
    attribute INIT_26 of inst : label is "4D2B336C8118F258250CAD46705402BB0F87C0C1F0FC7E631E0FCC60F60222E0";
    attribute INIT_27 of inst : label is "FFFF5577777557F557F7D577D7FD7FFF1D3A0B78058EF502190410C3C04000DB";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FB8A3A8081CDC93F10043C2446A";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "A480EAC280DD640080263924B2C96C90016CC01FD80C27E6497BCD6603636BD0";
    attribute INIT_01 of inst : label is "6400615610D5FA3944364C9B2D5143EAAE9FE14B6405A52B5A83597D393D67CB";
    attribute INIT_02 of inst : label is "4D17E8104A28E0228F0030ABD7299E420C06530CCA6306532F8402F90722A5BC";
    attribute INIT_03 of inst : label is "B2405B74058EE5E27ABFA001216C64CDF89FC6B81224A3F3C8000735662AF04E";
    attribute INIT_04 of inst : label is "862D9050B4EE2C0110AC013DB6644885AC7A8B16F01A855B41300868DB9A0050";
    attribute INIT_05 of inst : label is "27164A2D02D76622DDF04E00E8001D59845DB2BCF268AA84B405055500A28A46";
    attribute INIT_06 of inst : label is "D59785D26AE04788D4B56DA2404D14D84DB68A05D51B2A1C599832ED0657840D";
    attribute INIT_07 of inst : label is "BCF36A71645925D189B25DF04E05549680E63A814A0907F80E07E52FFD2C85D2";
    attribute INIT_08 of inst : label is "B7297DE27F4BA7BBC2D03362683C97B8AB2156E1C8F734BB0E012039C02796AC";
    attribute INIT_09 of inst : label is "AA92C6EB2C7E0B90F0D2B6E47AD45F5AA8A07BF426FD0DB5EC1FEBF9E9EB8164";
    attribute INIT_0A of inst : label is "677385ECA40002F651392CA91EB695AAB080ABF1CC523BA6B6A542C70F12AA86";
    attribute INIT_0B of inst : label is "0110004E100004400178452A93EFDF7274A04C435AEFA3FDFBE8D83F23F9F52F";
    attribute INIT_0C of inst : label is "9C9AC883DF781CA74802204C592B3B8D08965A0B3DA11653A2CF3BA4ACED9D00";
    attribute INIT_0D of inst : label is "B2D16C424CB2C2F9743200208BD5200208BD51CDDE3C50AB0847462A6BAF4F86";
    attribute INIT_0E of inst : label is "44C9AF142AFDB95E9092E6ADB6D171464910BD23F63D222DBBD3471E9252B6CC";
    attribute INIT_0F of inst : label is "A25E7A18C8B6EF4D84E3D240E50C617622A90540542E880054BFC5E32E4800E2";
    attribute INIT_10 of inst : label is "4079F3A31100F05522FE0064D0B3F9FBB42622A8008215188AA00208557377A8";
    attribute INIT_11 of inst : label is "22142FAF7A81F03E9A108252FC968284E221388B65689FFFB23B8204CDA10E08";
    attribute INIT_12 of inst : label is "74E3D4AA85CB57AF6A75CCB9484621A294FB3FC49B48C45D293DAA90CC435B72";
    attribute INIT_13 of inst : label is "AD6AB1595634D7658A36EE5A41483AAF7296C140EA00F25CCEDB69D8BF234D5B";
    attribute INIT_14 of inst : label is "D64F4A47B407F14A00EA0D4CCD98952880403F8E50CC8C480499006E2D07A96D";
    attribute INIT_15 of inst : label is "7749CD6F415538D55B5979DEFD290DDFFF7F1F8C4D485BD6D5509EAC2D69BBDA";
    attribute INIT_16 of inst : label is "461B9533BB15566118A0ED258769665E6DAF5DEDCA7A9EACFC7FC9B79C3DADBC";
    attribute INIT_17 of inst : label is "6127DE6B54B02F2111622CF3A39DC6F9927B114471B108ADBD9A78897672504C";
    attribute INIT_18 of inst : label is "20C8C9495CEF7295C3CF3CCC919B9CC5A0524A48C359E64ECE36A5ED636329E4";
    attribute INIT_19 of inst : label is "0D3BFF3FD0CB26221B2CC186ADBCE6CB1F2CD86E143A20CE234E14E840D83BB2";
    attribute INIT_1A of inst : label is "DE315720857211C628E40572123098668D1EC45551F17EA8FE54AE4292845E7D";
    attribute INIT_1B of inst : label is "86B2FBB044C04B6521E525B26FAA2DABF044555118CFF3C233887A498B61A3E0";
    attribute INIT_1C of inst : label is "BD1B208FC9B8A3874345821EE4A5CA72BC944788F3929C992E583FF7F64B6E20";
    attribute INIT_1D of inst : label is "000000179019FFC0081FF7E0381F80003802E56092E19EA7AB1C8F7F5BD6DEF7";
    attribute INIT_1E of inst : label is "6927D9BB89B337B6C9B9B9B9B55553553554CC00000000000000041111455555";
    attribute INIT_1F of inst : label is "8F0D10FFB4E483B6DAE1DDAE599F0B7ADC5705C1775C000E1AB031B418B09B96";
    attribute INIT_20 of inst : label is "2E7FABFE6B29492BAA31158CB50011231AD81F92081FCFAA8970964EDE2396BA";
    attribute INIT_21 of inst : label is "25D1BF1163D31C8D3FE8C4DA502AA03CA2482FD080031E85CF2273FC807FC440";
    attribute INIT_22 of inst : label is "3FE7B024000000200C5AEA35702094126A4C777DF00C462525C84E101B680214";
    attribute INIT_23 of inst : label is "EFB23F601ADD7A07DE4B905482E2492D83A280DFF56291882FFE2DFB995C6DD9";
    attribute INIT_24 of inst : label is "76F3D52B1F49CED9BD12C07FCEC0809E0000B0000782012A441C7C0D1D9E21A1";
    attribute INIT_25 of inst : label is "FC6E46E9377AB8CB2B48105C11AC8CC01157FE5BC4008BA12FC5132A536FBFCD";
    attribute INIT_26 of inst : label is "D96C997E3613D7332760FBD53B1B22F718CC60C3198C186333030E6031DABC6B";
    attribute INIT_27 of inst : label is "FFFF5577337557DFFDFDFFDFDDFDFFFF15F47D0F23EF7F2B576D79DA65660069";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7B970B8B8D8B90A67734C6D17F62D";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "B6D02A0085B16A1BA59A10000002090400207FD6984D37E548794D7719690A82";
    attribute INIT_01 of inst : label is "62680570D0025A10402486004930C06B44554158A6C4438230F5085D1E2F01C0";
    attribute INIT_02 of inst : label is "91016801061827128E3402B831D646800743AC87540D43AC870269BD44982128";
    attribute INIT_03 of inst : label is "8C6C1017A40B156051A2A0000834B00DB89D5408FBF683FB3A1A0004A7855407";
    attribute INIT_04 of inst : label is "81204C382523E90221E9020484400021A0518604AA0395C3444868000B1A2EAA";
    attribute INIT_05 of inst : label is "C10C3994C294A7809054070328DA05400709A2F85028EBFA86C4195501659386";
    attribute INIT_06 of inst : label is "1314F514508867A0A700FFEDBFF6E925B6C9759710820A00300A04081A813D10";
    attribute INIT_07 of inst : label is "A7945010C330C521E120505407057F50D8202A82D281C01D0250A9AB7BA8F514";
    attribute INIT_08 of inst : label is "550C050244382FF903065AFA030801BD3A8BC6F1C4F5140AC810384AE83CA098";
    attribute INIT_09 of inst : label is "A05AA4A1AA4A87E4F14551FAE8E8522923A3A1534850D142881FE1DF51720047";
    attribute INIT_0A of inst : label is "66414DB7B0D466DBD90DB8B6D9DB36BA71110B40D0921820A42092824F00382F";
    attribute INIT_0B of inst : label is "23F148EA22148FC523E88D0498B009823690BD0A023FB2401006903F297F446F";
    attribute INIT_0C of inst : label is "5EC2E80BF7557691297204666DBDAEE48C9FE66FBF66DF5D9BEB8EF6F6B7F485";
    attribute INIT_0D of inst : label is "A2CFB77F68A2C7817B599FB37BFF99FB373FFDB77B824C9BBDF6B3B3733BCFE4";
    attribute INIT_0E of inst : label is "616EF0932648D1906CFAFFE8A8897BF339B8F591DBA8DAAAC21A05DFDB2C1448";
    attribute INIT_0F of inst : label is "CE6051AD6AAB08689CB3FB71F2CE7B837B36D67E5E2B666FB7C3FE18AF4DDED2";
    attribute INIT_10 of inst : label is "665973DDDDA8DBC799EF3E74ECDFFF7E1B83FB367ECDFF8FECD9FB37FF6DDEF3";
    attribute INIT_11 of inst : label is "BBD770F36C85613E8ABEF77716A96C86D3E1B4FDB7ADCBFFDFBBC3336A31CF37";
    attribute INIT_12 of inst : label is "7A120A50052497F092DE1DAD2936050A52245004C38466617FB6C2526C0A1B7E";
    attribute INIT_13 of inst : label is "08413C9B8A690A14CFA2AF7145006AE97BD5C508F4C2B069F081400A69520156";
    attribute INIT_14 of inst : label is "868ED684207CA374475E4B42FFCCD4A4A8A3E51FA22FA66A66F8235A4B1B4E05";
    attribute INIT_15 of inst : label is "D0950B68C4A7AD8152124891A75AA4915A3762EAA8D552148051E486C1F8C210";
    attribute INIT_16 of inst : label is "2241052BAC524B25A8D5A9052B69449541484CA8AA51830F0821F10400214834";
    attribute INIT_17 of inst : label is "B145140330A048FAB22324BBA5DC263504135550110841297512B500543935FA";
    attribute INIT_18 of inst : label is "E040524A40E0708156AA2AC4808F58046011462C809064AAC324A9694145086A";
    attribute INIT_19 of inst : label is "4DF2AA2A127DB6864DF6C11429A820C84722D02207198A47BB02066002551AFF";
    attribute INIT_1A of inst : label is "A50637605AF618A0D6EC5AF61190C873E715C02370C168A0DF54B0F69A64CB21";
    attribute INIT_1B of inst : label is "E07A97A03BB00009002101242FBA39BE711023704E03F0C6112212008260004C";
    attribute INIT_1C of inst : label is "190A209551B86387D3C40002A455C5D15C2645D8B980CC0F43B8046120004E28";
    attribute INIT_1D of inst : label is "000000002A19FFC3E05FFFE3C05F9F03C044210084C80DA1286C018843188C63";
    attribute INIT_1E of inst : label is "880639CB37BC3871C1C1C1C1CAAAA9E81E843C00000000000000041111455555";
    attribute INIT_1F of inst : label is "06091F2AAEA44D245222090E53952EB3AC4E1384EF38013560A2C0A160A11C73";
    attribute INIT_20 of inst : label is "3EFFAAFE0A0B6D4AAB11A442A142D23AFA8C5D68433FB82AA452047FDE3B8438";
    attribute INIT_21 of inst : label is "0C8209051241A3A20660C1E05A83E84145142FE4E902222D592053D4A875C650";
    attribute INIT_22 of inst : label is "0AA7E80000000074DC91AD255A44A05B4A6C0CFF5068C1C12511461E124E2A55";
    attribute INIT_23 of inst : label is "83603C4003ACE258E843C93C49FC908B9AD5DF0888A0810C2B410DF0285A2D29";
    attribute INIT_24 of inst : label is "A20E150A0F50D1DA5A24C9AFF18000840004600023020008869E368ACC24CAB2";
    attribute INIT_25 of inst : label is "28AB61AC234AAA90837A804C737DFDCFD747FC5BCA9F8BAEAFC57A341A2597CF";
    attribute INIT_26 of inst : label is "DD7C029B8393B580334252903A162AA818CC00C3198C186301830F601C92EACF";
    attribute INIT_27 of inst : label is "FFF75DFBBBBDD75FFDFDFFDFDDDDFFFF1A3A295E37CBF42AC00D69DA25400069";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7E1E4BF84582850A5A7C742835628";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "924488E0854024AF76D20822820820D4410C542BD42B4DF9497E64D6D87889E0";
    attribute INIT_01 of inst : label is "28225067448048026804948001A280505444505B0FC60A0210940140252C200A";
    attribute INIT_02 of inst : label is "404920A0545101400211283330FA62041511F4D5084C11F4C10825A410512800";
    attribute INIT_03 of inst : label is "B0FE105308C95960C19284080331314484F5B8CEE9D241EF30A8A82601255529";
    attribute INIT_04 of inst : label is "014668A0042A6D0120ED01029F260441451D14203895419D0102A24020081C01";
    attribute INIT_05 of inst : label is "8828AD5686D201240055291B2088911D0241014040205000BFC4085F8430C282";
    attribute INIT_06 of inst : label is "1A1249E21AC2EA009C2EB6DB6DB65B6697EDBEFA0811A820A12A12080C681042";
    attribute INIT_07 of inst : label is "92231A828BA2848848059855291A0017FC045A0852A4420C5074A125482649E3";
    attribute INIT_08 of inst : label is "5F2295750A65221CA54F5ABEDD8E1C9E11EA0263A96E3DC9F454880A629118D0";
    attribute INIT_09 of inst : label is "28407241272CB76540C55D9AB06973AD3B49A87EF81D9866E60DF182713D5047";
    attribute INIT_0A of inst : label is "CEAB57B239F06BD9DB649C926ACBC234C1124A794A98296C9DB23508D400546A";
    attribute INIT_0B of inst : label is "62C318B823318B0C62A08F708A139894873DD00A63279B0310B62C1F132A6890";
    attribute INIT_0C of inst : label is "46C22A217757F73473FC07332CACCC69F74DBB2696724D08C9A1FE32B332F9CC";
    attribute INIT_0D of inst : label is "AA66DBA9AAA27315198C89113709C89113F09872738A9D3EC721919157D8E7C3";
    attribute INIT_0E of inst : label is "D16C62A74F4AD88726489ED1049D189996CF6B9D098E4CC6CECA59B86F2764AC";
    attribute INIT_0F of inst : label is "95A51CC6331B3B294A3F0DF6B2631491191262B747233234AE55924C83066430";
    attribute INIT_10 of inst : label is "234D22CC88A25CC9CD3313D2A64C062E49D119122444C9C664489113271C9CE5";
    attribute INIT_11 of inst : label is "CB6692304C6A804085CA592922EDB6C6D0D1A07EFA9E4E04CCB8F11923188B12";
    attribute INIT_12 of inst : label is "B254E808028016120262524E73B80538C724D6806D8022296190DCE7300AF84D";
    attribute INIT_13 of inst : label is "69CC0E13626F9B9044826501454262652857CD4812B5702AD7955E0962027148";
    attribute INIT_14 of inst : label is "9916042DA74283247523441212C4418E383A141D23212224D2C83A2764473A55";
    attribute INIT_15 of inst : label is "9890A443136C8B695A48AA95AC1036944053AE2439814ED69A6C42D524C8DEF2";
    attribute INIT_16 of inst : label is "239B39A8314862B4645D4C0CD3AB32120C3526A2A09D0B16682528EA20652947";
    attribute INIT_17 of inst : label is "412DB300B090820B2566360810503644821D451118084E2549D685E1984FA796";
    attribute INIT_18 of inst : label is "E14C48C101E7129D00B30FC718812A836A1168B6054C60AA6304EF2D3103CC23";
    attribute INIT_19 of inst : label is "48FBFF0E77AD9806F7B30414A54E309987922890255D8F4D591024622528435D";
    attribute INIT_1A of inst : label is "CDA3A6828CA811B464D00CA8198144B0601D615240C1693C5E308228CCDF6A34";
    attribute INIT_1B of inst : label is "766AE6383FE400010129A80001103B2470D95A400DC2F8A8A3023068D590206A";
    attribute INIT_1C of inst : label is "0A61E1413886404A0205041220D8CD0342A514B294D4A0D6F32C8C6900020922";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000010A9401145401003D6AB5ED6BD8421";
    attribute INIT_1E of inst : label is "F77802003FBFC0082E0E0E0E000002002003FC00000000000000041111455555";
    attribute INIT_1F of inst : label is "C050150BC5B455044200091D85760E338C0601806718050080E100E080E19FF7";
    attribute INIT_20 of inst : label is "2B67E4794124AD7352B1B9A91942D3B183B871A6413FCA82991A847B8C919210";
    attribute INIT_21 of inst : label is "00A3844E6711B0AD83144BD24CE02924D34D042F504414942A8F03D8C966A16A";
    attribute INIT_22 of inst : label is "233301000000019EB722A104327131C9555A4CFD3050B37589DC258B88029A19";
    attribute INIT_23 of inst : label is "8B046C401B8C6620C8B3051428E002088808A2228210940A333E0428863D9CBD";
    attribute INIT_24 of inst : label is "AA5AD439AF1A9B7B53FD680FFD8000040000204001000018059E15980E6E4080";
    attribute INIT_25 of inst : label is "CE01C1082A908E4980B0B1203E5F1CE25390BF3133D3E90DEBD11AB6147557A1";
    attribute INIT_26 of inst : label is "6C531BC1831660E151046F401802445A18C7C0C318FC187F01830FE05E80EDAC";
    attribute INIT_27 of inst : label is "FFF74CFBBBBCC75FFDFDFFDFDFDDFFFF19170E522BDE772192588C1880320070";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF86A85FB9A42880650E2274C067A39";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "2490381AA55504A6D36A132CBA936DD8518E95528C83C01351796C444D6D71E9";
    attribute INIT_01 of inst : label is "804813E09021701340125A2DA5451011414050412035146B5AA2452061B06419";
    attribute INIT_02 of inst : label is "690DC00908A28A02082409F0100011811A40001AD40340000C004AAB4059AED8";
    attribute INIT_03 of inst : label is "1200D92480B10F2E44B6120001800F4C049190A31224C30F1A12001406876830";
    attribute INIT_04 of inst : label is "0385514594A4CE05004E0516910C4885061A28BB62074F82042A5811B9101644";
    attribute INIT_05 of inst : label is "14514AA5146206876968302F61D2070045058330724051011000183F81A68A84";
    attribute INIT_06 of inst : label is "9462B0C618C8BC111B074DA69B49B4984892012497C2241145B48C2812E46D01";
    attribute INIT_07 of inst : label is "1507184515451885A2D609683028222203F101014B04093108E2C5442145A086";
    attribute INIT_08 of inst : label is "A4204A224858B5B0021E6B94C24D30082035103595E479B120208129886A34A3";
    attribute INIT_09 of inst : label is "019FC089F40891FF8707E41F403C8010AC80807E401B942C02981D0127600156";
    attribute INIT_0A of inst : label is "F6001636B3F2CB1B9A6DB2D6FCC9C63041112A6B1E5463CD18C05E017820A8B4";
    attribute INIT_0B of inst : label is "E40F390022F3903CE4008A629E32A99BC617A08C52A84F40226AC430554126B4";
    attribute INIT_0C of inst : label is "970AFD7C802A86182FA845767DCDACC0B3999E6CB1A6D9669B2C3B3736B7D0BC";
    attribute INIT_0D of inst : label is "EFCFFF03FBEF5B119B19BB77ED1D9BB77ED1982675060C15AC60B77731FBEC6A";
    attribute INIT_0E of inst : label is "EB705183046AD9C26DD8B2E1051399F33C9A5BED598CDA52D47451A8EBCD78FF";
    attribute INIT_0F of inst : label is "0D66198C694B51D13A351D68FCC635973776CEE156AB66EDC26BC65AA90CCC11";
    attribute INIT_10 of inst : label is "EE79AEDFBBD799E59A6376B26FD81E0C1B47B776EDDF999CDDDBB77E7609DD43";
    attribute INIT_11 of inst : label is "261CB2B3ECB80080D61983CB37BFFF44C411313FDA9CC400DC04C373E1F1BB7E";
    attribute INIT_12 of inst : label is "BA70D10004085A330BC66E8C2FE8462842A39227DDA26665A5D2C05F908C5C5A";
    attribute INIT_13 of inst : label is "318998D7CDF93054CDB3411C49090DC088A2C90A369CB42AD5128892A944458A";
    attribute INIT_14 of inst : label is "12A6D6A8C5B002F05A01A04AB6CCD084198D801382AB666BC6CA2C01A054760A";
    attribute INIT_15 of inst : label is "D370016300E060C58C5200529D5A14522180282A91D18C63114F3608D082D463";
    attribute INIT_16 of inst : label is "6475B038399144B9A08E0888A42A24A2082044C8EA1A294640360D2000463175";
    attribute INIT_17 of inst : label is "1539A2033111011BC64B28D0169126A59651186451BB5884E08A74A92266D368";
    attribute INIT_18 of inst : label is "2849924AD2E9153640E38D58311948066053706404016664CB32C72E2312CE27";
    attribute INIT_19 of inst : label is "498000846FC49845FA930C18C50C42A948388028969E8A4AA908976002040A02";
    attribute INIT_1A of inst : label is "E8BB1492EE49039770906C480BD8681A7408A751C8C16838E122B3EED8774CBC";
    attribute INIT_1B of inst : label is "D70AE0B833A42DB501A5AEDB6698127D71C751C9EFFC0F3022F6306D7B91BF62";
    attribute INIT_1C of inst : label is "7DDFE5753982F0810300419A40E02E0B8094B686F01280D9A3947FED924B2D08";
    attribute INIT_1D of inst : label is "000000000000000000000000000000000002C510144C6DDB70E6873DEE7BFDFF";
    attribute INIT_1E of inst : label is "0040020B00400000000000000000000000000300000000000000041111455555";
    attribute INIT_1F of inst : label is "4A080833D03CC8148A00CD4F256621C873D8F63D8060048B120625051205E004";
    attribute INIT_20 of inst : label is "40C04400210DE021FF1410A4124480A0853001A6101FC022A052956EC1851330";
    attribute INIT_21 of inst : label is "8AB3DC01A7041B8FD900081642720F2CB2CB102655211094A8A4801BF30611F7";
    attribute INIT_22 of inst : label is "0AB748004000838B04026515002212DC450195041244E8D29098B756D24E0900";
    attribute INIT_23 of inst : label is "2D9051FB18718E45D20AD4F2A79CD9FD018820A0A226DF131434402A2D5F67B7";
    attribute INIT_24 of inst : label is "2A423471708F08590324645F03F3819F9C0CFCC067E6033AD000581711960821";
    attribute INIT_25 of inst : label is "CC11F29EC83992410840B0E4D76B2F549D1A00A035648C71302B56F6D04E7811";
    attribute INIT_26 of inst : label is "06530E8101002CD83A035402380A0C5218C060C3198C186301830DE050D0CC58";
    attribute INIT_27 of inst : label is "F77744ABFFA847715FFBD9BBDBFDBFFF131B0DAA2A080701922DA88823200031";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF029C4BC3EC6CC12AC2B6C8A866231";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "B6D24C5A9B546640412911A69A4924DC0626FA52A9570A0DE17E82666BEB6189";
    attribute INIT_01 of inst : label is "A4E92042F24B285145924E6DA5410144540144499025040EF2872D2320112509";
    attribute INIT_02 of inst : label is "012CA1172820802432F49021492490924F4A490F5CC54A490965EA254C0DA6D1";
    attribute INIT_03 of inst : label is "9900C93794AD0531245A00000126202025B894A9DBB6980ABA5A44944B933C08";
    attribute INIT_04 of inst : label is "3365104094A607409207489090856A9525CA081B524801090CA96925B068C144";
    attribute INIT_05 of inst : label is "041042210C424B936B3C0808B27A49889F2D4C412B614410900008AA80A68A8B";
    attribute INIT_06 of inst : label is "8402FCF7C949260633242000490000490012490414CAC050409E01293AA43529";
    attribute INIT_07 of inst : label is "1752C94104410096E6D2CB3C08428012023348114B82837D282265C42144ECB6";
    attribute INIT_08 of inst : label is "ED6C4C224868A096103639B44A0C141D34AF0877A5683881F0B05229E9389420";
    attribute INIT_09 of inst : label is "0C68690E8690D244C0181092E3015118AB8D992ECA4FB32250C215423DBC2B57";
    attribute INIT_0A of inst : label is "0F0436A62480CB53D6292B948012442C03612931485329471090F23BCC45FDEE";
    attribute INIT_0B of inst : label is "08090200EC9020240803B62292020810A404203050806B197668408071123480";
    attribute INIT_0C of inst : label is "808A4A280A0234000820997669A988D044181E6C25A6D8429B097BA6A6269024";
    attribute INIT_0D of inst : label is "AA0925C85BEE3217D21112225511112225D116144A4E8549284822222DAD401E";
    attribute INIT_0E of inst : label is "524803A1522AC9364A94409B6F1FD1222C121D0510A4938288C071688208388A";
    attribute INIT_0F of inst : label is "490749084E0A2301D62D104AA08424122224944164B244493480105222488902";
    attribute INIT_10 of inst : label is "4428AE91112A51011202242648900A691202A224488951088891222545851292";
    attribute INIT_11 of inst : label is "2A5483ACEAA20C109D129248219248D494B5252024A884029486822253A13A24";
    attribute INIT_12 of inst : label is "B9365024941052020A40424808008828088696EC150044452110881041105C21";
    attribute INIT_13 of inst : label is "6118A05546AB0940892073452D0DAA711A67AD0FA351F8AA92371A9A8548550A";
    attribute INIT_14 of inst : label is "12A75E9185500F2095075068368CD0840A0A80790482444A148C4A877068265C";
    attribute INIT_15 of inst : label is "00CA50191FE3E88D185B0CD3B57A64D2611424AEF3D388C6135C2C1D82AAC8C6";
    attribute INIT_16 of inst : label is "6641301811534EB565450830B46426C6DB61846C6B4A07D7249301E0CE8C63A2";
    attribute INIT_17 of inst : label is "3728C636B2120C54078C24647368DE54925B28A22C994AA4C48A54A9AA520800";
    attribute INIT_18 of inst : label is "E749DB6B9DEEB634E869044D9199DC5C6453526C4A0892664592852422921866";
    attribute INIT_19 of inst : label is "5012AA045001201A0024102084856AA96822A16816B8964BBF2816E44A4496FF";
    attribute INIT_1A of inst : label is "A0B6AE86D8E86216D5D0DAE86BBA5D366CB5CD6B42C16822217C828C08264EA4";
    attribute INIT_1B of inst : label is "156E56922AB32DB564A7A6DB5110627F72256B42120D096BAA08036DC204D350";
    attribute INIT_1C of inst : label is "810C324A0C02D4522A2C934A6681281A129572AE5552AAD082B934ACBB692869";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000026724D5E8DF97E10E900421000010";
    attribute INIT_1E of inst : label is "0080040040000000100000000FFFF60060000000000000000000041111455555";
    attribute INIT_1F of inst : label is "082A7F2181862D14DEFB654E0162200803C0F03C000000000204040402070008";
    attribute INIT_20 of inst : label is "26886E84695B7129AADA158D955D0C44C039E8CDB4DFFFFD5EA7B57DC365B6A3";
    attribute INIT_21 of inst : label is "3EC4A8714A1A14B0A42A0C33E32A00E38E389C3FD51A774EF3D6900FF31251F4";
    attribute INIT_22 of inst : label is "B541D4000024034A4D321495132494105C1577043D994EE424B556765B68DA6D";
    attribute INIT_23 of inst : label is "0100004300000600C0020012008000180075D77DFD66F12A5C756E1BB85A2657";
    attribute INIT_24 of inst : label is "6E73952130D95E5BC17FC00C018381841C0C20C06106030A0000300000040000";
    attribute INIT_25 of inst : label is "04E3450D8800BEDA8941904533FD48C9035481E8A949A0E3601DE6F256C6C83A";
    attribute INIT_26 of inst : label is "D456388B3374B593F70AD020584BAC7018C660C3198C186333030CE00855C729";
    attribute INIT_27 of inst : label is "FFFFCCAAFEA8CFFBFFFBFBFFFBBFBFFF022A247AA25102890A2DCD99252600EB";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0652ABFF6C2C8DB22032F0AA52E61";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "002020307F45629964B238000000000400C03FF560472201687F46E2C97990B8";
    attribute INIT_01 of inst : label is "0110010100005008210000000061801451110508A27D8600041148010C010100";
    attribute INIT_02 of inst : label is "060140840C30C10B2C0800806D92D820908325D0A95A8325D60013A281200008";
    attribute INIT_03 of inst : label is "88261200086F6430F2B2000003111004A6CD693700000116442420029000440B";
    attribute INIT_04 of inst : label is "0001986100004100004100068F620440C0530C001C020406003080000D548850";
    attribute INIT_05 of inst : label is "861863318020900000440B182044040400008A2050001401824002AA84104044";
    attribute INIT_06 of inst : label is "C62000000070A0050800B24B2592DB2D92D92592CC900018612212000136020D";
    attribute INIT_07 of inst : label is "0020006186618820000000440B0280304E2430080080C0120C10808084030000";
    attribute INIT_08 of inst : label is "A7060217061415B1831308D001618629836510A3986700100C50180090C10631";
    attribute INIT_09 of inst : label is "08EAC708AC608BCC010002B200011884188385426D5098062C8A115E0363188E";
    attribute INIT_0A of inst : label is "BEE1A736B890C39B180DB0B6D2DB16B2C1520550808A10000846100040080020";
    attribute INIT_0B of inst : label is "20890820A3908224208288100C90688A17BCB02C18E86700002E7810755E0C34";
    attribute INIT_0C of inst : label is "C65020282220B7B7799807336D8DAC4D88D95F2CA9B259D6CB3A793636B6DDE4";
    attribute INIT_0D of inst : label is "C6A5B6797182838BD98CC9196159CC9196159966632078B0E625911111B9C42E";
    attribute INIT_0E of inst : label is "4364C81E2D008081245A5CC00003D89198D859B1592A4E2CC40C0D8ACB664144";
    attribute INIT_0F of inst : label is "242054C638B3103009B15974B66310811112722CF67B332DE6D6B20B830664BB";
    attribute INIT_10 of inst : label is "334506C88882DC9DCB3B931A245A0D4D89719113246599C4444C9196665998C9";
    attribute INIT_11 of inst : label is "FBF610B2AC61885035DE7B21135B6EC441F1106DB72EC282DF96F19968189B92";
    attribute INIT_12 of inst : label is "3000180003860A90C15228AF79981617F6E0D02499A02220A9D4C6F3302C352D";
    attribute INIT_13 of inst : label is "10842E01602998704586FB06B40B2ACFD804340831F0384091008404E0842080";
    attribute INIT_14 of inst : label is "09162108431E0B6D70E50C4E36C44DEE4838F05B6AE3622642CC38650C451282";
    attribute INIT_15 of inst : label is "09C18C00101FF2A09404E2040884A2040224A2A900240425082CC4402520C421";
    attribute INIT_16 of inst : label is "89CA0080870820300024040840AA1120001C3202028302060020601E20421082";
    attribute INIT_17 of inst : label is "43412142D5040F87F80FB2A8750D0E89248D4D354922942119508942008B6CB6";
    attribute INIT_18 of inst : label is "204428684062310C4010A8102A2B2A84AA841A9683D52489682448AA14C43168";
    attribute INIT_19 of inst : label is "02E95522332DB81665B7045842AA1008808C18CC207B0140410C21E205785300";
    attribute INIT_1A of inst : label is "3610C180435800420A304158009048122406840D00C169A4407EE1425EE22025";
    attribute INIT_1B of inst : label is "61901980445440001800000026CC0FF9F03C0D0000490A6211004E0052900218";
    attribute INIT_1C of inst : label is "134AF7D5088C2081010000001C350350D020540A81840C02C850A00100000610";
    attribute INIT_1D of inst : label is "00000000000000000000000000000000001000038854401000B40214A5294A42";
    attribute INIT_1E of inst : label is "00000000400000001000000000000FFFFFF80000000000000000041111455555";
    attribute INIT_1F of inst : label is "810C00927E5650810400482EDD251FF7FC3F0FC3FFFFFFFFFDFBFBFBFDFA0000";
    attribute INIT_20 of inst : label is "24A87EC710E04D10A87988000D724633E1080D16C97FE222BC5088EA8B318200";
    attribute INIT_21 of inst : label is "08CA880704058102800449DA8E240130C34D68002AD49E81A7A3D015F01570FC";
    attribute INIT_22 of inst : label is "ABA2C8004024911A18000820F011015A04071D843840D980080006DC48060000";
    attribute INIT_23 of inst : label is "FAFFFEBCFFFFF5FEBFF1FF8DFC7FFFD7FE00A82A0030708A386B055888AA3513";
    attribute INIT_24 of inst : label is "C618CF1080C0433838023FE8FD7C7E6BE3F35F3F9AF9FCD5FFFF8FFFFFEBFFFF";
    attribute INIT_25 of inst : label is "4A2B638484080001956221CC49259D32449140F2E34302E1C40D58208034C01D";
    attribute INIT_26 of inst : label is "2C26194B8300F580900629403000280918C3C3F318FC7E631E0FCC606E9089C0";
    attribute INIT_27 of inst : label is "FFFDC89EEED88DFBFFFBFBBBFBBBBFFF0C4CAB28234D0408130593F8CC100021";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8219CB890600866009B4481014230";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "802921387F04729B6CB42C924924924D48F27FE560450206667E0391C8789491";
    attribute INIT_01 of inst : label is "3014810909249D0C30492524906180105154055CA6458621083D0C8184419124";
    attribute INIT_02 of inst : label is "0C9274C08C30C3824B8A40842CB6584824A16CE4AA4AA16CE5D01340A36A124C";
    attribute INIT_03 of inst : label is "CA67B6904E6260369620000003353C43228A2E1E00002004C525304304489C49";
    attribute INIT_04 of inst : label is "683198634212531840531846CA33265070630C491D220427A214849349991A00";
    attribute INIT_05 of inst : label is "8618633181290449249C49D8040524264090922499341014C64000AA871C60C6";
    attribute INIT_06 of inst : label is "C629061C6474A6094B91964B65B2DB2DB2596CB24C904118624E22940116828D";
    attribute INIT_07 of inst : label is "483C646186618A411248649C49C20298CE25184C2188748A8C3930908412061C";
    attribute INIT_08 of inst : label is "02D7269523161520C391C6C12330C260816021830842823406710E845481E631";
    attribute INIT_09 of inst : label is "1A6883188821988CC120162264034CCE18114584256109930582015381419E8C";
    attribute INIT_0A of inst : label is "B4B1A4129C904209088498A24A491290CD928594218B84104A47326CCC1A6E66";
    attribute INIT_0B of inst : label is "208908213B9082242084E8980EB8EDCA533C904D18C82234DD0C2A00E5538C34";
    attribute INIT_0C of inst : label is "C2702A808282333679B8373324C4A459CCCB4F25E8B24BD2C96A3993129249E4";
    attribute INIT_0D of inst : label is "C6A4922B20828941498CC919214CCC919214C86321301838E621911111108024";
    attribute INIT_0E of inst : label is "49245C060F80A099244B584C3041489199C8CC914B324E2E651D048A5926D355";
    attribute INIT_0F of inst : label is "647264C638B9947408914B20926311C11112622C52293324B255170B0186643B";
    attribute INIT_10 of inst : label is "33C702488882CCBCCB09931C244E04448931911324648CC4444C91923218C859";
    attribute INIT_11 of inst : label is "CB6638118460905139CAD9638749260E22838884922670824AC271992C188992";
    attribute INIT_12 of inst : label is "2483188202C30AB8615728A679B83694E6D859249C802230ACD664F3306D25AD";
    attribute INIT_13 of inst : label is "94A62F01B230CC60448C8A823C1B1884540C3C1899F09B00A949A64CC0A530A0";
    attribute INIT_14 of inst : label is "4914214A530A1A4770A1048C124449CE487850D23AC12226464DB821048C95A6";
    attribute INIT_15 of inst : label is "8CC0860C30000230B504B3084085230884A4D0D10428252D4C34C0642838A529";
    attribute INIT_16 of inst : label is "9BCA90C7470C32300464804A50DA91286196132304E310049049201B325294A2";
    attribute INIT_17 of inst : label is "61C229D0CD400FE7FFF037A86D4B0D9B6D8EC71DC366B6330F718B66898924B3";
    attribute INIT_18 of inst : label is "10676E66705A2D6C211CB034EEE233819B8C8B9BA1772D9B796C58BA9C4C2158";
    attribute INIT_19 of inst : label is "8CCD55F133249826649304DA52B3380CA0840C8C60514160628C6153056A51A2";
    attribute INIT_1A of inst : label is "1690C512431108D218A24311088844302092650408C1694021C7B94274E23225";
    attribute INIT_1B of inst : label is "7193194844546490DA109249378D2D70EC1D04080219064388004B24D0910608";
    attribute INIT_1C of inst : label is "3342F750087630C32126482136352358D2606C0D814C1A46C84CE21249248534";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000193092C8964010049A46B18C6318C6";
    attribute INIT_1E of inst : label is "0000000040000000100000000000000000000000000000000000041111455555";
    attribute INIT_1F of inst : label is "B1849196005690C27186D82ADD0C000000000000000000000000000000020000";
    attribute INIT_20 of inst : label is "15881885DCA0059C0038CF18CCB2461161460A32C97FAA281C0068C883126A06";
    attribute INIT_21 of inst : label is "689280CF0634C3E28224338E1E20031861C76BC080770E08CF039C24B118785D";
    attribute INIT_22 of inst : label is "A100E0000100013A30186260AE9DCD4E880708803A4ED9AC6E0346DC480186C7";
    attribute INIT_23 of inst : label is "040001B800000801000C00600300003001AA002AAA9C30051C4BD196E82A1513";
    attribute INIT_24 of inst : label is "8318CF94C0F4733E74008013FE70001B8000DC0006E000300000400010100000";
    attribute INIT_25 of inst : label is "5B9A6D84040861B6A52441884805BD36C4B180C2A74600E0800E48298338B018";
    attribute INIT_26 of inst : label is "B484D94262204D0633B67BC1B5A029090000000000000000000000006FB199C0";
    attribute INIT_27 of inst : label is "FFFFEABFEFFAAFFBFFFBFBFFFBFBBFFF0CEEB3002245881C21833114C49C0084";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF909CB0A2020B6600BA60A11185B4";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
