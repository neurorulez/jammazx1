-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "4BFFD0783552C0EA03129A75E6E9AD84B7FFD4FFFFA9FD793DFCC581FDE7E7DD";
    attribute INIT_01 of inst : label is "04A2191115D54BD8B09FFFFE585E76517DBD5B895A92EB013445FB7B96A1E59D";
    attribute INIT_02 of inst : label is "FFFF6FFBACFFF88BD608AFA84AD121DDF85C81427792B8A2A86C3091996452A0";
    attribute INIT_03 of inst : label is "CE7FFF151F8387F17E481A09068240D0481A0906827FC12EE919274257FD98F3";
    attribute INIT_04 of inst : label is "3C7C4F9F7A39E0E1C5BEB63AC32037F1E77BFFFE1C151F8381EF602000203038";
    attribute INIT_05 of inst : label is "B6B6BFF829837FD01C83643FFF97F466001F07FFE1CE1FFFBFFFEE73A75C11C0";
    attribute INIT_06 of inst : label is "5DDDBBBF7FFF545319C2E0181D33817CEDFE38BD7471A7E3DDF9A87B394AFDFF";
    attribute INIT_07 of inst : label is "0E7DD356BE1F5EBC3CF9FFFF3610D26203F1E9B43F1FBE7CCDDDFB32D590601C";
    attribute INIT_08 of inst : label is "79FE78FAE7A9ED3FDDFABEF351F47FC1FFFF2C6839E3EEF5C3CB55D952846020";
    attribute INIT_09 of inst : label is "FAE000DFF736F05F2E458326DC7CCB780E6233EFA7DFFFF002410DBDF667C62E";
    attribute INIT_0A of inst : label is "BC7FFF4955690479F77BFA91037CC9FE49F626233332161DF3D1D7B7FFF48212";
    attribute INIT_0B of inst : label is "7F92678DBADE9BBFFFEA8A8FEC5154CD29F7A40237FC1CE1CDB8FFCF80DAB68F";
    attribute INIT_0C of inst : label is "1743F3F6362B33951595257DEEFFFFAAAAA8E9CDE27B334DC9EE58028FF14032";
    attribute INIT_0D of inst : label is "890B26C9B3ECF8679E57FDE298F53C0270834FD37951416D1DA1AC1F2E6AE32D";
    attribute INIT_0E of inst : label is "39FA6EB52AA7F66A0891046073BFAF1F90C44FD360C0DFEF39DFD27EFA4929A9";
    attribute INIT_0F of inst : label is "06FD3FC4622CD7F900F7FE403527EE2FF86273AAB67FFE98FAFDC05C81DE7BFF";
    attribute INIT_10 of inst : label is "6ABD268D4783490429F0173FB00D76E8841CDA6936ACB595CD26BE18830DE000";
    attribute INIT_11 of inst : label is "18C9ED34E69A53CA6BAA9ED3CA693454F0D375442CE9A27CA947DF6880997ADA";
    attribute INIT_12 of inst : label is "C8C8B4D8CA873AE62478F1E2D88E66D8A5F34C594A688A9AE648462305B4B44C";
    attribute INIT_13 of inst : label is "9F2CD193237DC60C8FAE79CFFC85595B8C66B718D18952E304F6C7D590886B6A";
    attribute INIT_14 of inst : label is "63FFEB1C7DFB7A4231414C5216E919B24492C9B3C957DF6FBEDF7DBF368D122C";
    attribute INIT_15 of inst : label is "25DF393F8B4E33642CE69FBB6C803BFB3FF47E3600802B492CA54B2C4544DFFD";
    attribute INIT_16 of inst : label is "700005B88A960618AA635C4588F6308C9EAEDF4ADE90BFAAEC62BACB4AC9B274";
    attribute INIT_17 of inst : label is "BE4804EADAB6CDA362D723E8F7DADB211057A12ABB7EF2211F59D519B3C9F9BF";
    attribute INIT_18 of inst : label is "06F3E491B23A71B2DE493E69AC4D34CD345336600B0C5D2C86F991576DA018EF";
    attribute INIT_19 of inst : label is "FECFEDFBE5B1FA5559A0A4E52A4C6BF79AA5F3548FD8B20000000F24FBB00054";
    attribute INIT_1A of inst : label is "ADB671C924E28F96ECE4058370EBECF96700CECE6CFA5BF7FFBF6EABCF5A7A77";
    attribute INIT_1B of inst : label is "8583D91A11B860229FCFF664CB2532C942C79FD1E843045E40C5E0091C6D1A36";
    attribute INIT_1C of inst : label is "4AD4FE1BEFBFCB2F2C02D81591B759ACE001AEE4F3B4425EA6E58AF58A666EAA";
    attribute INIT_1D of inst : label is "AA34B617EF8A0A2C27CF514FAE8EF24EBC9E57FA9DF01709FFFFFFDAFB6DB6DA";
    attribute INIT_1E of inst : label is "E44748550B0029580150B00A88A5601515C731047CDAF37E75C36A1696C9A406";
    attribute INIT_1F of inst : label is "DAB5A727CDFBDE406B6339068542A7FE5D3027DB694A8AA1441010BB7FB37327";
    attribute INIT_20 of inst : label is "ACF3BAF05498FC0A86992798E39B2DD7FC7E02E7A9ED9F4868F64F2018F6F5A7";
    attribute INIT_21 of inst : label is "57D60C8262A55B6DC49E5AFE6C8E9F245E48B058186E2BAAB4D96A88A6227FAA";
    attribute INIT_22 of inst : label is "98857D2664BB5324B4402CF93FC4200C7F659806AFB6B930BC925E12CD0C59A2";
    attribute INIT_23 of inst : label is "92AB43F2EBA018000600202026606575B1DF2783FD8E792F35E4BF27063E5576";
    attribute INIT_24 of inst : label is "0100505400050404FFFFFFFF23F7A068A965760BC55CCBCCBCE9406D2A349416";
    attribute INIT_25 of inst : label is "A95DDFFAAFEAAAAAAAEEFFD57F5555552A9541D4F50493940198000066404000";
    attribute INIT_26 of inst : label is "3C0000000012586C905B6000C00AA01FE060600000111117FFEAB5553FFF55AA";
    attribute INIT_27 of inst : label is "044444444441111111111110411192A000000F5AFFFFFFC200010115B6C9268F";
    attribute INIT_28 of inst : label is "BB98A5C10E2170498A8C42CD4000000004208000108003FF9102244089111111";
    attribute INIT_29 of inst : label is "2236414422235505A2AA211046AA08B451518823BDEEF7928C4A31BDEEF3BBBB";
    attribute INIT_2A of inst : label is "145520822254118A2A9040018A08C50548208AD504668AA4104566A235455088";
    attribute INIT_2B of inst : label is "508352120809482118A112A410404A1108C509120908094046282A410404A823";
    attribute INIT_2C of inst : label is "D3D9FFB3D23E93778EDCE94B7167FF778E07BB9FDFE3EFD3BC59F350FFC9808C";
    attribute INIT_2D of inst : label is "BEB97F9B7BBBAEA4ED70CDC3E5F1C3CE067267CC34B3B258384E6C5F478EE1F4";
    attribute INIT_2E of inst : label is "6369D7527BE6A7301A7CD8FCF96359FEBD4D2649F96DBD68CAC68CC040EBC37F";
    attribute INIT_2F of inst : label is "003FBDF6FFF6B3447CD9199DE4CF62EBEF3F1B42BA97635BC1ADE36D6749E7DF";
    attribute INIT_30 of inst : label is "954AA000000000C444D1BABAEB105BBB56ED7B5C288A70DF4EA8089E00000000";
    attribute INIT_31 of inst : label is "A1B4569715376982D2E2A6EECEE5A5C54F7CB75ED3859996BBBA6B9599A5552A";
    attribute INIT_32 of inst : label is "95444FF7711B5444AA2211BFEEEAA2211B3686D3D3CE9E3686D24F49E3686D0D";
    attribute INIT_33 of inst : label is "33333811EAAAAAAB335C669A69A6AC14F7A9999999666666F299990626663E5A";
    attribute INIT_34 of inst : label is "B6D2355556AA5555555884D2764435557DF95DDFDF8947777774C0777372064B";
    attribute INIT_35 of inst : label is "26405E826017A3542767CFFF1176ECA4103D36621AE93FD51CB5FFFFFF773721";
    attribute INIT_36 of inst : label is "65C9D6E14BCD0D3B2D12FF10DB34A6D4DB191D9A58F06A542774202EB7D79017";
    attribute INIT_37 of inst : label is "4ACF520444D93B49B2626AB934AEDBAF34D4918C3F5E474C9CACE9D6C174D9B7";
    attribute INIT_38 of inst : label is "8570947568A334D3E7066BB66A4440D1774E2018524A494929A536A4D4D29352";
    attribute INIT_39 of inst : label is "80EEC0B97C2BE14B026500240000AA65C5A549B59F2D0AF27C608D9AF3F3E6AF";
    attribute INIT_3A of inst : label is "D61475AE031D77125C0C312389A412ACC92E63232777633B9A69A73E80FE80EE";
    attribute INIT_3B of inst : label is "26008841C313862C53882E15E0370AF00AAB94154ED4543B5154ED5FE802A634";
    attribute INIT_3C of inst : label is "AFF97BA63673739CF4E67FD6FF9FFFFFF3F77703127511345AABFCF155555150";
    attribute INIT_3D of inst : label is "5867B54F9E222FEC135434D7FCD82774D9C1B019C01E7F3EFEFF3F1FF7F7F27F";
    attribute INIT_3E of inst : label is "1EE18010200202B9FF7FC4EE57205C76D1180A81DD2C3DC76D5274C65C365DAE";
    attribute INIT_3F of inst : label is "FF9CAED9B41292FCF7EDF2E9D21690EA364F39F532F52DFFDFD1CB5F48D7F8FF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "D48009907FF7F968B386397F8C60B569980091BFFEF3C793FAFC8B13FC0EC79C";
    attribute INIT_01 of inst : label is "F6E652832A8A818C340008FECCBCA46FE9A28D19AB8FB189EABC876CA79E8A97";
    attribute INIT_02 of inst : label is "FFFEEAA0A355521EB5A1EBFA9FCB68448EF82A9F48B4C3E8061129B3DDED7ADA";
    attribute INIT_03 of inst : label is "F5CE7230854AE623016AD369B6DB569B4ADB6DB4DA6001F85CB53F8BBA321BDC";
    attribute INIT_04 of inst : label is "E1FF372775C71F1E3E3E46E4FD9DC69EC55E10860130854AE0631CCF3F9FEFD7";
    attribute INIT_05 of inst : label is "80011293842D6ADFD7FC9FFDB71365D9BFFAFBD5FCA36A52E4A421084318E567";
    attribute INIT_06 of inst : label is "2DD65446CCCC4000D6796EEFEDEC7F3BFE5686CA4A9E1D9CA23D462EEF398969";
    attribute INIT_07 of inst : label is "77FEEB575D479AADF317A72B0003A39C7DAFE453EAE795AA229564CC49DE5EFF";
    attribute INIT_08 of inst : label is "76EB2FD4CAAFB58D655A4EA88E559EBFAD7B0003A63DCE79A8D7552A5CFFDFDF";
    attribute INIT_09 of inst : label is "FB5FFB2FF7489F9B2B1A72DAEBB78B7FF11DF2B19935BA30003EF25EF792BFAD";
    attribute INIT_0A of inst : label is "FAD5B4C000ADD5ECF85BBD2E7D8F74BF3256DABDDDDFEBFAF9DFD75D54EC200C";
    attribute INIT_0B of inst : label is "3FCCB4B6B962CBEAAE2040628A956576EFF74BFCDFFFE65EEDDEFFF4FFE9DAE2";
    attribute INIT_0C of inst : label is "F775D979B6F399AD6476D4939DA56980014A2AED7DA4DD9EF4EF2BFCE7FA7FD5";
    attribute INIT_0D of inst : label is "54C481304191619003E542016D12C19F6117506008001D95EEBDDFECEFA9298A";
    attribute INIT_0E of inst : label is "0A0C01DAC44D5A93DDB8599B001606404D08D06016097530800D2C83C59474E4";
    attribute INIT_0F of inst : label is "00647FE57B5477F88A27FF329A0D8CF5FB14342ECAC7F96501818C9693000AA1";
    attribute INIT_10 of inst : label is "800A56609FB983A157EC66C1D7B6205C2F3BCF18EDC5ECB8781365C7D564E000";
    attribute INIT_11 of inst : label is "99C098122FF6C12026B40981A0346098034A98AAF50E1AA976B42966E524F9AD";
    attribute INIT_12 of inst : label is "AB9D564B9F5D4DB99DEB57A97A56FA9950068DBBDDE524195882A9152ECA12B2";
    attribute INIT_13 of inst : label is "68D362249DB338F795DFAEF5470C888671B70CE30A37619D7A870F2605D3B68D";
    attribute INIT_14 of inst : label is "0E6DB071C46CD1B9C2CFB4ED3B1E656D8BAE2A40B26A05940B281640CA52615B";
    attribute INIT_15 of inst : label is "DE28C6C514AAAA4BE2EAE88D902AC4955FE923564B513C36DB7F069B88896492";
    attribute INIT_16 of inst : label is "122226CA31D4DCA31EAE6A895B956A3B2D36E0371305F01D95944CF335B56DAA";
    attribute INIT_17 of inst : label is "6182B72D640D369D876DE577440F640BA48F9004C0A23E0ACDB2266240B20611";
    attribute INIT_18 of inst : label is "6B28385E55029AC623E283DBFEDFED7B7F0DEFD65D5EAB5EFF96A59924847310";
    attribute INIT_19 of inst : label is "0130B2042A562CF9AB45DA2F72E4A4AD0BD88A8D100108CC899912584F8B549A";
    attribute INIT_1A of inst : label is "4001428002A5A86980EB3954D7121334B5BA8B5F902F2C81040993FE30040499";
    attribute INIT_1B of inst : label is "0A962CD1CA4184B440001100DD6EA55A85701B12DFEDBEDC33EDDB71E62DD916";
    attribute INIT_1C of inst : label is "DF4B9EE0B2045D50D002E95C2004069159989141D232153E5EDB71F2908B3175";
    attribute INIT_1D of inst : label is "00A13222D1D465F50A22F7CA4BC3808B8008002F470C81F4FFFFFF59FDB6DB66";
    attribute INIT_1E of inst : label is "588882B66DCF132E6D265CDB72C9B9F2BD79F3DA24598116A251283F5D42C668";
    attribute INIT_1F of inst : label is "47334A825624003BFAC640F6488D020102CA504D95937E4CBA6FDD00A08CA829";
    attribute INIT_20 of inst : label is "50480FE3F86ABF9514E22AA8C319210423E1900A92B941EF9551550BA604BB70";
    attribute INIT_21 of inst : label is "8B19BB34A7C6800132E60139711122C7E597D7AF27D17C75F204911134441455";
    attribute INIT_22 of inst : label is "B99C9EC60533D55BF2800BA608088115D0AADCCCF0CB46C7CB7165EF3C93F590";
    attribute INIT_23 of inst : label is "772C8EAC288CAB534632A242467D05895768C31C8AA30232D65ECBE6DC8A3C95";
    attribute INIT_24 of inst : label is "0440010001100001FFFFFFE81D80C4B3501294BF9B415CB5CB4B8CB3725AB8D9";
    attribute INIT_25 of inst : label is "FC00000005555555404455557FFFFFFF0884634A10800119990BFF0077111110";
    attribute INIT_26 of inst : label is "C0000002EC145041105043FD40154015587F980000ABABA000001FFF955555FF";
    attribute INIT_27 of inst : label is "441555400511005004555149051483E0000002AEFFFFFFD40001F150209967F0";
    attribute INIT_28 of inst : label is "547E02F01FA8FC07E80D2976A00015AD45010400000FFFFFC448811220154441";
    attribute INIT_29 of inst : label is "EC203226ECEBE6991193B74624649BA8C8DFE6C2B7EAFFEF56EFFE6A55845050";
    attribute INIT_2A of inst : label is "C969CE4EC2225D64B4E72661112EB24A7B93B08C97512D3DC9D844CBAC969E64";
    attribute INIT_2B of inst : label is "24A29CC93B088A2DD6494139C9D844416EB24A9CE43B08897592539C9D8444BA";
    attribute INIT_2C of inst : label is "2423C010500135002B7802987A0800002AA962AEE07DD40406820331FFC412EB";
    attribute INIT_2D of inst : label is "CDC38035FBE393DAB60AA80A583D7A42C0014801D546006D760C36E010400E1B";
    attribute INIT_2E of inst : label is "C58549EC265BCE1C7D986E9733BCE51A4FB6D5752EF66AA5F7BA5FFAAA3DD9F9";
    attribute INIT_2F of inst : label is "00037C42B60A4589586E55535AA9AF7CBF12E4064F6C85A052D0058495989072";
    attribute INIT_30 of inst : label is "198CC552A954AA5050C5045145FEEBEB5416EB56ED7B0C79C670DF4E00000000";
    attribute INIT_31 of inst : label is "AFF5F63FDC7FF5F6C7FB87FF6EAD8FF707DEFF540019011A3323B22A221A6633";
    attribute INIT_32 of inst : label is "B4451F77DC714451A228C71EEFBA228C71FEBFD75ABFFFFEBFD76AED5FEBFD7F";
    attribute INIT_33 of inst : label is "A5A5A8BCF3333337018A4A28A28B85615FB12D2D2D787878E6E1E30661E79F7B";
    attribute INIT_34 of inst : label is "A69373333398CCCCCCC8D2460985900028A9088A8A8007FBFBFAE0FBBFFA66ED";
    attribute INIT_35 of inst : label is "5102B295062C2EE9F48B10135A8D147497F042AEA0A018072084FFFFFFBBFF9B";
    attribute INIT_36 of inst : label is "AE156A1A26B86CC540EFFF5D445000000153442803F766E9F4830EFC67A052AC";
    attribute INIT_37 of inst : label is "01EF2FFFD12B88E2571C651050000A5E48CDDABD8012D805F5C501797E014280";
    attribute INIT_38 of inst : label is "2C064B7A400E500C35130001E6EB02FC58A90BDF04A082140010000201282085";
    attribute INIT_39 of inst : label is "3E88160B03421A00502C00050000C1A8D6002F32B1B2740CA192D619C5858670";
    attribute INIT_3A of inst : label is "504CB330312CD23160480314012427060C5154445101100005B649C13E093E19";
    attribute INIT_3B of inst : label is "2A00444A090412032020702C33181619818DA203560C0D58303160DDC0207113";
    attribute INIT_3C of inst : label is "C8285248A4A46529554800B8A80FFFFFC6545502635130224145143117151150";
    attribute INIT_3D of inst : label is "5A822B9E00688FE723F73754154909232D863F75FDF0040200A8801510065282";
    attribute INIT_3E of inst : label is "E1180210000017E3FCC3D719201723168E64AD3E8040C03168A7833C80F41190";
    attribute INIT_3F of inst : label is "C405F0808A29260501103F122CA121CCC87500D2462F60FE401DBF8999300200";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "32280482CAA518219A84280A6A6510690ABF917FFE539283F9FE8301F80FD3AC";
    attribute INIT_01 of inst : label is "E0E6028102A280CC0407F4028C0000AE8D064195910D219DC4B8142EB506C180";
    attribute INIT_02 of inst : label is "FFFFA5522EAA9BC4E6BC4F7A854748C8EEA2AB55512082403A0113A595B95090";
    attribute INIT_03 of inst : label is "55B9CE648A8FA3E7FE0AC160B259564B2AC160B0581F8CA25DC08BCBA947D015";
    attribute INIT_04 of inst : label is "D085D44C18DA6F6ED88888541D6FC116E739CE725C248A8FAD8C6E479FCFC7D7";
    attribute INIT_05 of inst : label is "F6B62D69888C1507E97CA9D64D44908ADFE4F92A4CC66DAD9FFF7EF7855C628B";
    attribute INIT_06 of inst : label is "C08C95593FFEF4536A9E06E3EC8DBED524AA1B9470A6AA5D4CEA8B715A5278FD";
    attribute INIT_07 of inst : label is "F294855412490630CD66FFFBB61140AC3D4E1883D56AAEB45CCC995410A76EE5";
    attribute INIT_08 of inst : label is "CA141B28212A4512C8AA90510EA0A95EFFFBAC69DACD2A9049005400043B8FCF";
    attribute INIT_09 of inst : label is "022FFB49B41267941008754A0D890753F62CC1411AAFFFB8025E7494A0A158CA";
    attribute INIT_0A of inst : label is "04BFFEE9550B6C90202040063D01505410A0484C4444E2E410465583FFE69214";
    attribute INIT_0B of inst : label is "040428109102889FFF3AAAA504920410520841FC4091E82E900B00103F0902A5";
    attribute INIT_0C of inst : label is "62582081E2410101242048A00273FCEAAA0840108C814500500009FCA0025FD0";
    attribute INIT_0D of inst : label is "47570BC2F13C49E486B2A6E38D770D3F51965FE11D514F21600E01E84AA94004";
    attribute INIT_0E of inst : label is "7BFC2210000519D3A2AD59D54008254EEA8CDFE10B1B51562040F0FF0E37C757";
    attribute INIT_0F of inst : label is "03F76A85F36C4D50CBEEAA32DA0F68F7FB9237CF0AED538D62AD489E93521153";
    attribute INIT_10 of inst : label is "CFF7E414C5096BB55142643155151556AE30C71C7D4768A9AD4A7D288D54E000";
    attribute INIT_11 of inst : label is "7C4A0141120854128096A494129004CC71BBECCCDCEB9AE9FCA532406DFC50BF";
    attribute INIT_12 of inst : label is "E35D77C35DDA6ECC42952B51B4DC4CA1236AE82BD543B9907EEAFD172F6E66CC";
    attribute INIT_13 of inst : label is "3597FB3FEFE9CC5D5B50DF1A5FDB3B33D9D067B3DBBAF0E62EF7DF9755FEF1C6";
    attribute INIT_14 of inst : label is "CD3EDE6DA5B670D162CAD8E62E6B34B70D54EB375B2DBADFF7F6EB6DF0DC3B66";
    attribute INIT_15 of inst : label is "88B5839734E4996D4ECD36FEDAAEE7DD75503E787211BE7B8621404ECCCFE7DB";
    attribute INIT_16 of inst : label is "E32326FBB1F492B39EE97C8D9A6673A5BE3AFB19CDD5ED86D9F76E9A0664B70C";
    attribute INIT_17 of inst : label is "0FEAE7ACB6639E1725EB56D7D71FB6AAF6C50006E2ABFCAAF96D7B33375B6B8D";
    attribute INIT_18 of inst : label is "7DB6D45B673AD77C56A85820348082A0909E84245610B0B51F1D7CDCDFE47FA6";
    attribute INIT_19 of inst : label is "9B3D5B6C2A577CEDBB75FD6F5AA8DB39B36D3AD5A951F79DDF399DEFB596A9CE";
    attribute INIT_1A of inst : label is "1FB7233F6E66A6FCCECF01D615ADB1BCD695ED57CDD534FEB376DD5579FA2FDE";
    attribute INIT_1B of inst : label is "DB163CE847F964BBA97BFD20077B11DEEDA2B0D0F08400232302F00906081014";
    attribute INIT_1C of inst : label is "9D8F56FC3CFAD75DF803515FC781F8FD79180C41F2A15714048198A0184086B1";
    attribute INIT_1D of inst : label is "553192E9DFB662B5E846B54525555E08843E14D58AA8F154FFFFFE10F1F8E074";
    attribute INIT_1E of inst : label is "4EDEEAA3478A1B3C513679A9A26CF353594F2134F8105F9EBB5F0E3D9D9BF32D";
    attribute INIT_1F of inst : label is "EA21667DBBD252150302AA440CEDA8DBC71EFFFEDCF9AA7CD4340A12AEBFE73D";
    attribute INIT_20 of inst : label is "029A651B2C2A291D9FBB3E1C92486190D5151E2E1985FE8FFBCF7CABF7F1E4AA";
    attribute INIT_21 of inst : label is "0DCF2597C776D827AEBCD1E75B80DD613AFA6930355A76B6A0C4D5B9B76EF180";
    attribute INIT_22 of inst : label is "611B6360E7CCB694A1C00053158CC91930AAD8CCFF6FEB5475C33AB8639B1D02";
    attribute INIT_23 of inst : label is "A9AEE9D763E8BA322522E3232441A0CDD5B56187CEAB379D73A8755492916B67";
    attribute INIT_24 of inst : label is "0001000110001110FFFFFFE508C7CDA19B52D6ABD52BA75A75E4D8DA9A6C4C9D";
    attribute INIT_25 of inst : label is "FC00000005555555404455557FFFFFFF773BB3D6F58082210908006644000001";
    attribute INIT_26 of inst : label is "E8000003E8268009A08203BA00176019807FE00000ABABA000001555155555FF";
    attribute INIT_27 of inst : label is "000000000000000000000000000083E000000001FFFFFFD40002015430C107BA";
    attribute INIT_28 of inst : label is "515EAAF55782BD55E281039940000000017ADA44000FFC001BA776E9DD400000";
    attribute INIT_29 of inst : label is "50208284505208A1141422828450142A0A15050D4A8500000042A54011295005";
    attribute INIT_2A of inst : label is "0A2105250B29210510828395341082984141408A08454420A0A0410420A21050";
    attribute INIT_2B of inst : label is "287A104414ACAD0A1050E420A0A5659A508286505314ACB08414C20A0A565042";
    attribute INIT_2C of inst : label is "B68BCC9198073D1526FC2BB53BBFCB1526AD4FF3B7A69A575EEFF211FFE46108";
    attribute INIT_2D of inst : label is "EF438437FBF2FDFE6F7A65C9EDF4E950DA172FE5414703DDFE7E2EBD5B52EA6D";
    attribute INIT_2E of inst : label is "8EFCFEFFDFED4F1A6FDC5E7E3B7F2C9FF7FDF364FD2D8CF868CF86BBAE1599FD";
    attribute INIT_2F of inst : label is "000ABC5EAA9FFECD3C5ECCCCEE656B7FFFEDB7E7F7FFCEFB877DCEFFF29F6DBF";
    attribute INIT_30 of inst : label is "1E0F00000000005500D5015015041045BAEFAB5416EB56BC3F0C79C600000000";
    attribute INIT_31 of inst : label is "FA9FCB4022804209680458000512D008B20900B632333230100011101000783C";
    attribute INIT_32 of inst : label is "1AFBAD7DD2010510D7DD011AFBA828820153EA7F76ABB553EA7FDAFB553EA7D4";
    attribute INIT_33 of inst : label is "0AA05B80FC03C03E5240679E79E6240AF051A8550280552A2200AA692AB01E68";
    attribute INIT_34 of inst : label is "B49530F00FAAFC03C03988447312177730635DDB0634E62266208E6AAEAADD2D";
    attribute INIT_35 of inst : label is "A21356AA33552AB555156BAB45124835552366EC8AA808B11694FFFFFEAAEAB9";
    attribute INIT_36 of inst : label is "EADD0CAA87AC68135949AA401004210421D2410208A043B5551D0A92556190D1";
    attribute INIT_37 of inst : label is "808A1AA545BAB38B7572414404210A316E8552B58B56DB457D797916EA22AD12";
    attribute INIT_38 of inst : label is "AA048269E9880474259A484342BD42AF5448AACA941290524849092124048010";
    attribute INIT_39 of inst : label is "BAA9570A1552AA8550280000000082AAD0000220B0857D3F54A62AD05A2AB416";
    attribute INIT_3A of inst : label is "0004A5891229623E120533E24086122448A2188108080808AE1B6EAABA2ABAAA";
    attribute INIT_3B of inst : label is "1A002881210242141342291DB0148ED81605122C144CB05132C144C82E058129";
    attribute INIT_3C of inst : label is "6BDC2D6E9AD656B5B5AC5CAC5E01FFFFF4F66601204101052ACADCD354411550";
    attribute INIT_3D of inst : label is "9381AA9C016EFD5E3AA71713ED812DB12C04825048D0209AB85EAE2BD5C1BAF2";
    attribute INIT_3E of inst : label is "B7188010410005C3592EB19FAAA737448728E2AE8540547448579FD416649500";
    attribute INIT_3F of inst : label is "CDB5FCCAAEB9B4776557BFDB70BDB976675C8AA3746B44FE4A19078BD1014251";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "07A82AF862218C9313AA3987BFEE4C628AB5737FFF9964D1BBFFC281FAA4F184";
    attribute INIT_01 of inst : label is "804260092A2AAA86624C17564AC630B5450AD0FEB4CEF2EEEDDD330887265340";
    attribute INIT_02 of inst : label is "FFFFA5587F2A88AC620AC438EDAF70CE84FAA7D394B9344069A0A9291A181012";
    attribute INIT_03 of inst : label is "2806300A35500803002008040000000000000000000007550886892F8B43CD50";
    attribute INIT_04 of inst : label is "071A0B33E624909123776783C28022A918C40002A24A3550027381B060301820";
    attribute INIT_05 of inst : label is "8948D2963563EAF814025209B23B6E25200A06D5B1291252400020003AA39D44";
    attribute INIT_06 of inst : label is "3F7362268000CBAC1541F818134240285355A42B8E515182B315748C84850000";
    attribute INIT_07 of inst : label is "0D2B7AAAED16F9CF1290000349EC1F53C2A0E5780A95514AA33366232F58900A";
    attribute INIT_08 of inst : label is "35EB6457DED4BAAD37556FAAE15F56A0000153942522D56FA2FDAB7FF3C03030";
    attribute INIT_09 of inst : label is "FDD000B64BED906BE97702B5927678AC09531EBAC5000037FD818B6B5E56A335";
    attribute INIT_0A of inst : label is "DA0000D6AA74132DD5DFBBF9C2DEADAB6F5FB7B3BBB91D0BEBB0AA78000D4DE3";
    attribute INIT_0B of inst : label is "7BDBD5EF6CF557400065150ABA6DFBCF8CB73E03BB6E16D16FB4BFCDC0747D4A";
    attribute INIT_0C of inst : label is "0DA7DB7C1D9EBAFADACDB656B500009554B6BFEF736EBAF5ADFF76034DB9A02F";
    attribute INIT_0D of inst : label is "554743C0F5BC69E58622A6BF852F0776FDD199691AAEA05E1DF1F6159554BBBB";
    attribute INIT_0E of inst : label is "932D2210000BADDBC5CD4C9A5008B72AED4E18691277BA532840F0C11E1D5545";
    attribute INIT_0F of inst : label is "07FD9558AF2A47FCF4CFFC287F85F4EC1BEA13E01E6FFF853B27CACD18D61953";
    attribute INIT_10 of inst : label is "E4997B6467D96B353CBEE3C8F37AA246AC8FE69C6C6676C9151072CCC5A4E000";
    attribute INIT_11 of inst : label is "2228D91A749B51A2365E8D91223604563CD754447E539CC388B87A7777FE2D72";
    attribute INIT_12 of inst : label is "5FDA6CA3D98EAB56683061CFA378BDE4B73CFEC8C677A3BD3D6A3DDF2766EBE9";
    attribute INIT_13 of inst : label is "7D17F15E9FEA977D8F087F0F378C7C7529E8EA578FBBD54BBDABCEF5D47BC742";
    attribute INIT_14 of inst : label is "5F924A78F31330D37EFAF987ED335DDE943053DB7D3C9AC935926B25E87855FD";
    attribute INIT_15 of inst : label is "42BD174352EEBB25056C7EAECEA62B6F3FE388A8725CFF7F5D6D56955557B249";
    attribute INIT_16 of inst : label is "43AA9EE13DBD9F935B6715CED3FBD7DFD31D3ABAD7D4CD4B59DEAB7FBBD5DE95";
    attribute INIT_17 of inst : label is "6BEA71DEB2FEB836BD8B63C3B1FBB3A9F562D02A3ACA97A8D4EDD591DB7D2F1D";
    attribute INIT_18 of inst : label is "659255096314F963662A8349BDCD26ED36DF274447893D199E957D47692D4DB5";
    attribute INIT_19 of inst : label is "8A3B592AE2F15BCD3AE52E6316304918912E14E1C3C0922B1F751D64916B3444";
    attribute INIT_1A of inst : label is "64937BC926D72EF5656CFC87D3EDABCDD2DE65C3F6D974268134C8477D6E1BFE";
    attribute INIT_1B of inst : label is "AF927A7CAFC9A67F2D4AAF62978365E0C79B9BABBCA2820BBB28BBCAAE07FD0F";
    attribute INIT_1C of inst : label is "B98DF279BAEA461DE2A93D3BC58A4A24B1CC4A30FC3B538B76FEACFB766EF6AA";
    attribute INIT_1D of inst : label is "55DBB823FBDF952C3A7636452464D3858C52146169AA9D24FFFFFF1DFFC0FC0D";
    attribute INIT_1E of inst : label is "A4756A33179718BCBE3B7871FC76F0E3FB4F7B1F4C1DD2AFDFC21B75918D62BD";
    attribute INIT_1F of inst : label is "85BAA636EFD8C626A5ADECBF4447A04B770E24DEC8CD9466CB768FDACAE2E14E";
    attribute INIT_20 of inst : label is "56D239898838968A9B919E3DF7DF7E9476B5539E2984DA9F7ECABCA8F6D576CA";
    attribute INIT_21 of inst : label is "94E55FDECE74DC24A63C72EABD81B7E09FD97CBE7498E6267AE3DAA8937AB1D5";
    attribute INIT_22 of inst : label is "254DA5E1BB889E5E7AC0127F946EF7FCF0E2AAA3F8672F4D3FC29EF8E13B09D3";
    attribute INIT_23 of inst : label is "88CEC77EC1A8B22B378A6E3736346354F2FDF29F479A6B0FF1EE3F2E8EB14DAB";
    attribute INIT_24 of inst : label is "400400884408C000FFFFFFFDD646FBD8A9C3F3154A1DA3FA3DB460D88C6D473D";
    attribute INIT_25 of inst : label is "FC00000005555555404455557FFFFFFF7FBFC10A40841101090BFF4288040444";
    attribute INIT_26 of inst : label is "4852852850144829104A210414A895401E7E0000CC54545000001555155555FF";
    attribute INIT_27 of inst : label is "0000000000000000000000000000815000000000FFFFFFF40004C3B830C10452";
    attribute INIT_28 of inst : label is "E919A0CD466833519BD2D7FFE0001EF7BB7BDEAF000000001FEFF7FBFEEC0000";
    attribute INIT_29 of inst : label is "45208A24114208890451208A241051222890144B9DBB7CADF2F56F953E53BEEE";
    attribute INIT_2A of inst : label is "82A941145208894154A08A290444A0AA5045148222505528228A4511282A9411";
    attribute INIT_2B of inst : label is "0A2294045148208894145128228A411444A0A294115148222505528228A41112";
    attribute INIT_2C of inst : label is "B78928A0683399B0AED4388F53FD6BB0AC0C49313486187074FF5FAFFFC0444A";
    attribute INIT_2D of inst : label is "9B1933927E8B252CED5CED7B2C75EBD26619672530D21A58784A2C3DCE938945";
    attribute INIT_2E of inst : label is "9BED92976DAE655772F458EDB96129DC925D07FDDB2D84CA984CA9AAEFA74C00";
    attribute INIT_2F of inst : label is "003E83716FC492C6745A19DC2EEF422E60B4DF7494BBCBECA5F45BE936CDB6AD";
    attribute INIT_30 of inst : label is "201000000000001111D5000555015015041445BAEFAB5406EF56BC3F00000000";
    attribute INIT_31 of inst : label is "012040A200020900144000449040288008200204001011001101111001108040";
    attribute INIT_32 of inst : label is "15005A802A115005A8028115005A80280124048081540A2404800500A2404809";
    attribute INIT_33 of inst : label is "550AAC08C03C03C2A404400000000680028102A855552A8022AB540020081990";
    attribute INIT_34 of inst : label is "8000300F008843C03C0680518400100040190004018007773330C47773322648";
    attribute INIT_35 of inst : label is "B209655B33D9963D39566AB83D9B6F22CAF5B6864FA89BDD3F8CFFFFFF773301";
    attribute INIT_36 of inst : label is "E36EBDBA875A5EDB6D90FF3C9926224449B023933C5A763D3954D1792288525D";
    attribute INIT_37 of inst : label is "24DFA55AB6F8D02DF1A9362326224145BEEC6A10CFF2DF746C7FFEB7E7A2CD9F";
    attribute INIT_38 of inst : label is "A81002E060052653495D8890F63F018DD675A9A911A226448891122244488911";
    attribute INIT_39 of inst : label is "A7ABD70DB752BA875036000100008CE60E01827B887F4D2B66DDECBD9BBB2F76";
    attribute INIT_3A of inst : label is "0C44E185123873300A112301422412E449BA22A2A22AA2318E1B2D4FA7ABA72B";
    attribute INIT_3B of inst : label is "0E001480A981532101A0250480128240080710101C4440711101C455CE021205";
    attribute INIT_3C of inst : label is "57D22D6D1AD61695A9AF5C8A5199FFFFA4B22404300202020CB8888220222260";
    attribute INIT_3D of inst : label is "BA7B4CCB8E323FEE362FDF8BE8B1CE6DB85F3469D3EA1106BA51AEAA25C1A4CA";
    attribute INIT_3E of inst : label is "F71800000000057936EFEF3C44B3B48FADB6DFB8B51A5708FAF61435A7F537DE";
    attribute INIT_3F of inst : label is "E890B9186CB4BA5C36571799F0BD9537329C98A96A6324FFCA3AFC2FAFA34151";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "94AAA8DC40A519DE5291168A0C990C6442A545BFFE5B1AC380FFAA5AFE6DDAA3";
    attribute INIT_01 of inst : label is "A2C142C2A82808E6C6069502A0AA0036885A8531AD4D7E89CBD804B315069A6A";
    attribute INIT_02 of inst : label is "FFFEB559C22A9C04E6C04CB8054844A8E4A02B0110A00140F0400DA25539A150";
    attribute INIT_03 of inst : label is "0011000008400283AA2841041041020820410410411550888002F92B8514110A";
    attribute INIT_04 of inst : label is "2423110004000000828020110C800C0002110826080012400002400005010080";
    attribute INIT_05 of inst : label is "812001205A1000808064510000050000808428000291C0201882601205003011";
    attribute INIT_06 of inst : label is "804004027248CA6000008544440D14400A0040900102101C084100602008A281";
    attribute INIT_07 of inst : label is "7402000092AC05000031948B4010044262020200B40002094104150000050D40";
    attribute INIT_08 of inst : label is "061880A52A810040900420440A23420002414280104402001421000202122222";
    attribute INIT_09 of inst : label is "8208A4000802258048881C500100035AC0886440101204B42506960400290100";
    attribute INIT_0A of inst : label is "45245848C02440934800000828081A0680801204984020A08414882485041841";
    attribute INIT_0B of inst : label is "82205810070A209098201112156600110C00400828802516800414CA24680015";
    attribute INIT_0C of inst : label is "010225110004450000B4A0C08A12808210914008C8822113323088205024D404";
    attribute INIT_0D of inst : label is "52425284A4A82900863AA4370D3E073487B959051A8204000144404A10C14558";
    attribute INIT_0E of inst : label is "9B20A2100000101BA2885D1400C850AE0A7D1805096D29520020E0C30C125242";
    attribute INIT_0F of inst : label is "0300003A9535A556EC5AA9FB5B4D43EA0D8C61E80EAD530724263D9914421552";
    attribute INIT_10 of inst : label is "6DB12055C81383A1560EE0F1415214442E23C69A6C5450CE1A0C40A90491E000";
    attribute INIT_11 of inst : label is "D570220D1B64A05418170620D40A99DCEBFDDDDEFBCF1BF9FDEF3804458481B2";
    attribute INIT_12 of inst : label is "D040786041C26F0CCC183165A95A1962C6FBE0CCC6443301ECC2A3973224D2F7";
    attribute INIT_13 of inst : label is "640D9730C6DE4C5C891E4BC9CD8E666C9CEED93D8B9937262F65CDC70543960F";
    attribute INIT_14 of inst : label is "0136C80C367BE7C5EE29F0AE3C4FC6EC8E69CF7F2D2DB84B7096E12C685AC179";
    attribute INIT_15 of inst : label is "5274164E5374DDFD9CDE6944482AE7FF75423070EF1AB51E59128150CCCC26D9";
    attribute INIT_16 of inst : label is "8E7357455528025550617FABF07F7F06DF3CF899CD857C46F8D66E323F96EC8F";
    attribute INIT_17 of inst : label is "0AC2B7AF12CC325E17A72245C661120A84CD1006E4AD670BC93F7F777F2D6312";
    attribute INIT_18 of inst : label is "64B6D0192732E360563269B67796D9B6C9C6489DF6633273381E05DDFFE6FFB0";
    attribute INIT_19 of inst : label is "181909626875608C3B6525631738DB39B32732F5C141B73B3E767C25B0F2ECCE";
    attribute INIT_1A of inst : label is "4DB7A39B6F67B6359CDC03CF959B81BCD696EDD2DFC0356E237049411ADC624A";
    attribute INIT_1B of inst : label is "8B38B8614869BD3DA142B0EDB763FDD8D58A87527184104C6704701D23018194";
    attribute INIT_1C of inst : label is "918C72B855C8A69C609A479B64D8DA6D7FAA50E9DA221520581A190290CBB449";
    attribute INIT_1D of inst : label is "0079980B5BD604CD08563DB56D444089CDFE214528888093FFFFFF81F0000004";
    attribute INIT_1E of inst : label is "4ECCC2FB97A1DDBD0AB97B199572F633395D2317F911403BFFD03921819DB22C";
    attribute INIT_1F of inst : label is "0BA2626D8990429DDBCCE0744CC5C34B161AFFA44AD58F6EC630CBD4AA0B673C";
    attribute INIT_20 of inst : label is "09B30561AC3A819997332E0E5971C1E15191102E188DB6AE49C65C0A8DB1DFBE";
    attribute INIT_21 of inst : label is "0F9505962470C041BCF811C658052C6158C2653335784606A200D199B7667020";
    attribute INIT_22 of inst : label is "03AFE5A0E7A2B696A219824BD118DBB822E82090D224231CB1C05838A21B1114";
    attribute INIT_23 of inst : label is "82C6C146877292EEA18B4EAEE00540CDF5B46187BFA0102C6586B3208281CFE7";
    attribute INIT_24 of inst : label is "989A26120241AA42FFFFFFE44DD576939842CE4CE6100B18B0D163D82CED162D";
    attribute INIT_25 of inst : label is "FC00000005555555404455557FFFFFFF7FBFC14850049201090BFF42332882AA";
    attribute INIT_26 of inst : label is "591A14890004000900020010042AA4C00079E0CC4855555000001555155555FF";
    attribute INIT_27 of inst : label is "8AAA2209A2242AA0AA2A0A868A8AA50500001000FFFFFFF400000338A2882116";
    attribute INIT_28 of inst : label is "541988CC46723311980848001B5BA2520100005000000000000000000104228A";
    attribute INIT_29 of inst : label is "5028A2851452AAA1451428A2851514228A114500481022142142044204214050";
    attribute INIT_2A of inst : label is "A2215145028A215110A8A2814510A888545140A28854442A28A051442A221514";
    attribute INIT_2B of inst : label is "88281505140A2A0A1510542A28A0514050A8821514140A28854442A28A051442";
    attribute INIT_2C of inst : label is "96E80AE69093B4902428944003414A90268D4BB3B4A6982888D05A21FFD0510A";
    attribute INIT_2D of inst : label is "2548F80204026D24433044C16CD4817866C120451937C80411044202A5754844";
    attribute INIT_2E of inst : label is "B250B692DB6D6DC66248845912101089B6480330B2030CE010CE011054571407";
    attribute INIT_2F of inst : label is "00114201940DB24D288508C86C6428C6C06D9285B496C259F12CD25372DB6D9B";
    attribute INIT_30 of inst : label is "00000FF8000000BEBEC0000000000000000000000000AAAAAA0002AA00000000";
    attribute INIT_31 of inst : label is "01606AA200A8DB4D54401845B55AA8803AAB68A842222222223332332330FF80";
    attribute INIT_32 of inst : label is "10000800043100008000421AAAA80006212C05800800402C0580200402C0580B";
    attribute INIT_33 of inst : label is "55000A10C03FFC035D0C7FFFFFFEC57FF831AAA800002AAA6254000420031492";
    attribute INIT_34 of inst : label is "49262000FC007FC003FD0C4A69C315DD80017FF80018C511111048511110224D";
    attribute INIT_35 of inst : label is "DA19B49DBAE92630111A73981ED9B244932E9BE48990BB66A36BFFFFFD111121";
    attribute INIT_36 of inst : label is "A3A139CA041A48EDF624AA99806141E83C024030A1A2463011102653C8710A69";
    attribute INIT_37 of inst : label is "D1003A64AA68EB94D1D344426149EA72988C67948136F1B45452113A42236ED9";
    attribute INIT_38 of inst : label is "2A4B6ABFE60861609C59D27B4621018C98E90AE4A0540883106A0D41A9152624";
    attribute INIT_39 of inst : label is "022997001952CA865000000120008184060036020C340429A490F6819DADA077";
    attribute INIT_3A of inst : label is "5E000234A100800E694E10E529C2620588DBB323333B33248C1B244A022A02AA";
    attribute INIT_3B of inst : label is "3100704A90152022204074A8033A5401912821224080890202240817C804403A";
    attribute INIT_3C of inst : label is "4E4BAE6FDCD75694A5A4118F48B3FFFF80000000000000000000000000000000";
    attribute INIT_3D of inst : label is "303922D899111D463E07D71B26110C49268ED8F6EAB66730234808E9011992C2";
    attribute INIT_3E of inst : label is "B9180000000005CB10A68710881538604C248E088606584604C25854D444C517";
    attribute INIT_3F of inst : label is "C9B513B92CB9B150295EA50961F89976665E48C3616213FEDC283579D5218761";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "D0DC82F1755759E85681976EA6637B60658E84FFFFA0BD0842FC8B13FD00D7AB";
    attribute INIT_01 of inst : label is "A1DE4A972A880AE7D41A78A834BE60A2A170141381AD346FC28907F72DA628BF";
    attribute INIT_02 of inst : label is "FFFF0FA0B47D58A6B60A68F2A718C3B1E5AF0300236249C0200447B3777D3050";
    attribute INIT_03 of inst : label is "1000042408400001992248000049124008012492001988A0A0A58DAB93983121";
    attribute INIT_04 of inst : label is "040220000C0001108080A01004010C0000012126000010000002020104000480";
    attribute INIT_05 of inst : label is "80008500521080882044100000411000840020020290C0A03804640000807010";
    attribute INIT_06 of inst : label is "041215021040C86008080500000C3040000040300902A2080041004028080289";
    attribute INIT_07 of inst : label is "4442001292A40500012080A32280404016020340340120094400011000054900";
    attribute INIT_08 of inst : label is "043A88A102200040101000051021420430410010086040001424420020811240";
    attribute INIT_09 of inst : label is "8281042008028504008938000108014C8080A844000240349100944401280900";
    attribute INIT_0A of inst : label is "2D21444A0804D2920820401821091A458080110408C02001065D020005041800";
    attribute INIT_0B of inst : label is "92600012051230108C320410872C10110804514A2000815CA000348200308011";
    attribute INIT_0C of inst : label is "A100351100415400001128800A1200A284012000C0AB00103210848451069480";
    attribute INIT_0D of inst : label is "1818641906C1B1180A77485201C419558D7DDA072D2284800140484211400450";
    attribute INIT_0E of inst : label is "2B40E41000045517999E0862811F18F319BB9D0724C1698CC0CF40A808101818";
    attribute INIT_0F of inst : label is "03052AAC85ED0553A6EAABBDDA61515C15FA3500001D5201C0DA0A9B56202BA4";
    attribute INIT_10 of inst : label is "DFFFFC4EC817313812057877C157EDCF2481C6986CE4C1980343E1999E8BE000";
    attribute INIT_11 of inst : label is "8A180F008924F00E03D780F01E0101CDE3B0EDDDDDDFDFED8005B48555C4D1FF";
    attribute INIT_12 of inst : label is "EC64728465A2660DDA142855A55948874A62D0A8CD0621616CF03156B8FF5AD2";
    attribute INIT_13 of inst : label is "8EED933886D80D59BC48E31D01AC20201AF04030AB5B7006ACEFA983606228A6";
    attribute INIT_14 of inst : label is "5176CA8A303374C56A28C2D6AE8B0481CC20DB371B2FF9FB71B6E3667D5F0562";
    attribute INIT_15 of inst : label is "E13EF0A75267996D0DCD2051FB0266DC35578069D2977098E2B7C220DCCE2ED9";
    attribute INIT_16 of inst : label is "BAEAEE1FDD642B75565530B815604755B75DBD7BBFE05EAFDAD66692262C81CE";
    attribute INIT_17 of inst : label is "BEF02DAD7E41455755D66F1180047EC0C4C8100660356EC0C61B3B77371B37E0";
    attribute INIT_18 of inst : label is "6DA6F43B66B6C3608E78149252B2499249A6DDB54EC776D7787544CCDB655DEA";
    attribute INIT_19 of inst : label is "4DDD1B350142E4BCFFEFFCF332689BBD376D36D5804125B8AF715C49BA8264CD";
    attribute INIT_1A of inst : label is "4DB73B9B6E57673E0DCC01D6619BDD9CDF92EF00CDCA366E1B73FEAB9ADA36C2";
    attribute INIT_1B of inst : label is "AB5D7A514C576DB412E76809B4076D01F504455679CA20A0EFCA729B2650B12C";
    attribute INIT_1C of inst : label is "D7BC403282D87FFE740909D93225F9FFF57B6C4C216381344808190255D99C19";
    attribute INIT_1D of inst : label is "FF2DE5FC9C96A4609D8E7CEF6E9EE9FB153670FA1DCACE0BFFFFFE81F0000006";
    attribute INIT_1E of inst : label is "4ECCF02BB7A3DDBD1CB17A35B366F46B6A840612DCB1E9DDBB09F9ADADBB6AAF";
    attribute INIT_1F of inst : label is "5962786DDB40028CF318732C4895E0BD2C026DA0DECD8F66C6B5A9203556C3ED";
    attribute INIT_20 of inst : label is "81BF8A955421E899973B6C6AAAAAA9F0F8F959EC1E0DB75ED986D8C0C5BAED9F";
    attribute INIT_21 of inst : label is "4DED4557156AD701ADB4A9A6DB0C4E633CE66732B75C571722BAD199B7666208";
    attribute INIT_22 of inst : label is "E77B7B616DD547132310B6E3903BC75A29816AB9C46C33F07980BCB1845A2315";
    attribute INIT_23 of inst : label is "91D6F167036ABEA6A82AE6AAA98C80CDC1BE7D87AE15565E6BCD7A28222CDB77";
    attribute INIT_24 of inst : label is "1A10269008490048FFFFFFEEE4F560B19AAAD66EF623479C79D8E2D91D6E8E2D";
    attribute INIT_25 of inst : label is "FC00000005555555404455557FFFFFFF7FBFE2DEF580000109080042FF822000";
    attribute INIT_26 of inst : label is "9112048BFC209040209042BC04354040187E18844855555000001555155555FF";
    attribute INIT_27 of inst : label is "108288218804822800808084100086A510541000FFFFFFC00000C00904124AA4";
    attribute INIT_28 of inst : label is "A91968C3465A30D197F2DFFFF430C0422B7BDEFF000000001FEFF7FBFFFA8A0A";
    attribute INIT_29 of inst : label is "0020A8041502AA01054020A804154022A011500B9F3E7CB97AF56ADD3A7AAAFF";
    attribute INIT_2A of inst : label is "02810150020A81014080A801054080A040540082A04050202A00415020281015";
    attribute INIT_2B of inst : label is "0A80100540082AA0101500202A0041550080A8101540082A04050202A0041502";
    attribute INIT_2C of inst : label is "04501C84330E0A00631020948A9B970062AB7BABAFE596C242A6EA25FFC05408";
    attribute INIT_2D of inst : label is "688187B2844E6F6C713444D16CF0E91B6211244D1500AE6061C83033295648A9";
    attribute INIT_2E of inst : label is "E6E4B7B6DB6E81EFF6D0605B21812491BADE12B0B7338CCB38CCB3FFAFA88A82";
    attribute INIT_2F of inst : label is "001B4260370DB6CD30624CCC6E458996D06FB73DBDB6F6D99B6CC6E363836DDB";
    attribute INIT_30 of inst : label is "C0000007FC0000BFEAC0000000000000000000000000000000AAAAAA00000000";
    attribute INIT_31 of inst : label is "FE9FFFF755FF6D97FEEAA2EEDFEFFDD54FFDBFDC62332233323322323320007F";
    attribute INIT_32 of inst : label is "15555AAAAE215555AAAAC31FFFFAAAAC21D3FA7FF7FFBFD3FA7FDFFBFD3FA7F4";
    attribute INIT_33 of inst : label is "AAFFF618FFC00006030C6492492584000071FFFD55557FFFE3FFFFDE3FFE1492";
    attribute INIT_34 of inst : label is "49262FFFFC44C03FFFFF0C6001CE1D550007D5500078840000000C400001040A";
    attribute INIT_35 of inst : label is "D405A99D4B6A6670023AB4D44EEDB06CB32CDAEE9D789F433021FFFFFC000021";
    attribute INIT_36 of inst : label is "373370C20E3858ED662CAAC982E1E95D0A0B4A70F1A3C670023804774D63336E";
    attribute INIT_37 of inst : label is "199A32748349E70693DAC5D8E1E056E2D18EF3BF99AEF5AEC4C0837240CF56ED";
    attribute INIT_38 of inst : label is "08224A60400CE1C13B7BB8164771029CB1DBC0E0708E13C07A4741E81C038470";
    attribute INIT_39 of inst : label is "004D04145841C20C1C51000000008185120067620E9401DDB8B27531ADCD4C7B";
    attribute INIT_3A of inst : label is "3F0808406002020080E000081C00220088DCAAA2AAA2AAA8080248520046004E";
    attribute INIT_3B of inst : label is "00FF008C00180000200440420220210100706200E1880386200E189DE8400200";
    attribute INIT_3C of inst : label is "CE495608ACA0E5294541939ECCF6FFFF80000000000000000000000000000000";
    attribute INIT_3D of inst : label is "30356104067A354EBB57B77D263549692D2CA09542908C0B26CCC9B9993696A2";
    attribute INIT_3E of inst : label is "9B0100000000074049F69358BBC1380C0E2CA6004B017880C0C0705409640916";
    attribute INIT_3F of inst : label is "DDBD44C86DB5B0F0E18EEC5B4039B77666DC88CB60E68BFE4C22115DC56D8761";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "83FF90FC6AA08CE813821D0376E0086087BFDAFFFFD17E9141FCE1E8F9C5F29E";
    attribute INIT_01 of inst : label is "84452048CAA00982404FFE56466C20E1C5D04C98900FB408A48490A7E71669AA";
    attribute INIT_02 of inst : label is "FFFEC550032A9B9CE6B9CC0F9DE366EC80F480409D3904801908A3A898288302";
    attribute INIT_03 of inst : label is "00000040201008A544489269A6924493429A49249A621822882C8A9F8EC59C5B";
    attribute INIT_04 of inst : label is "404000000011080800000000010A480001020802A8402010081010000048A102";
    attribute INIT_05 of inst : label is "8108200042180100008000220200004002210800021088080280200001400019";
    attribute INIT_06 of inst : label is "00400010000040800010010004C0010002125201012000000000021100002200";
    attribute INIT_07 of inst : label is "A900000004A02000084004010800000020105200000008210010100080100100";
    attribute INIT_08 of inst : label is "0000A01020000254420041040200009108030880000200001480000088044010";
    attribute INIT_09 of inst : label is "100004010008480012800920400084022080000000090C1000020020400C1040";
    attribute INIT_0A of inst : label is "114000C4124200024000010210000210800420020200002814008000220C0040";
    attribute INIT_0B of inst : label is "802410000040A204006040101100402020690820840001000040400090400014";
    attribute INIT_0C of inst : label is "0004044080044C012000100281402180001100011100080102408108124C0200";
    attribute INIT_0D of inst : label is "2121C2709CA72D62AE02BDF082E11C05B13E1F89D80800008000102800000440";
    attribute INIT_0E of inst : label is "73F13A1000011643C481085925A97BFDAC99DF89D14DC54F92D290FC12292121";
    attribute INIT_0F of inst : label is "7CBF556DD13A12ADCFED5773F6848C5C11879FE01A22AC82F63EF9DB1FCAB95E";
    attribute INIT_10 of inst : label is "C5B3672467C249040DF867ADD01C3340841EA28A342C24818510374E6126FEDB";
    attribute INIT_11 of inst : label is "0A48911264921122241689112224244420924644584310E9A0A4367045923CB6";
    attribute INIT_12 of inst : label is "EAC57382C596224731B366CC935CEC136124CE1960F0849C6C480416396C22C8";
    attribute INIT_13 of inst : label is "3B0DB11212DCC45D875B3B679D8C9099886333118B0B1A632C218DB19008C102";
    attribute INIT_14 of inst : label is "CBB6CE5979B360C16208D8862C13999684B243B65BADB2DB65B6CB7B60589165";
    attribute INIT_15 of inst : label is "45BB195616EC3B64242CB772DC8022DD0AAA5E2CCA5BB2DB45484484444496D9";
    attribute INIT_16 of inst : label is "E262673F1164177996CB1688D2E35F2DB70C361885901B02D8D623DF82519686";
    attribute INIT_17 of inst : label is "4EC801DDB7321816058761D59BB4B7201067C022362DEC2014DB9111B65BDB0E";
    attribute INIT_18 of inst : label is "6DB6DC0B6210D97266088A49084924C924B722405719B90884909046493459ED";
    attribute INIT_19 of inst : label is "F69E5BDAA2D036AEBD626E6582045B39916C90C9B540B7180E30196DB50B1044";
    attribute INIT_1A of inst : label is "249371C924C32DB4642C059611DB69DE46D8CD42ED9D936CFB66DD56DEDE26E4";
    attribute INIT_1B of inst : label is "8B3FB80C61337FF25FCFEF20076B01DAC59B3CE976B1CF1667317C60DB8E1C87";
    attribute INIT_1C of inst : label is "258ED231CF33F7DB6009BDFC8B12DA6E733C3E10E638409F37F48CF913366C98";
    attribute INIT_1D of inst : label is "00298820DE563394227613256D65B286B43611F5EB609136FFFFFEFCF0000009";
    attribute INIT_1E of inst : label is "A4444801C30C0E18611E30C0CA3C61818D167858D81CB2983342862DCDCB722C";
    attribute INIT_1F of inst : label is "8E382CAD9B2D423353039CC70445A1FE51052DB2D850B02859164CB62F76C90E";
    attribute INIT_20 of inst : label is "F5B9ED912D089708F6910C9C515145D1EF2C122C8B2DB68ED892192011B0CDE5";
    attribute INIT_21 of inst : label is "85842C966572C8258436C0B21D959B6496C9309810995656F8404888D66324DF";
    attribute INIT_22 of inst : label is "333B636421A29658F8509B3B2798C31977A2709CCF6C1B012D9216B2490859C6";
    attribute INIT_23 of inst : label is "8CC2CBB6DB70D8242643642026726445D1BB6992EE817B0B616C2F661636EB67";
    attribute INIT_24 of inst : label is "10128412A8610060FFFFFFFB5AD726E88B02F6F2F8DDB2DB2D766058CC2C6605";
    attribute INIT_25 of inst : label is "FC00000005555555404455557FFFFFFF1C0E104A10800001090BFF4203028800";
    attribute INIT_26 of inst : label is "1D1204895430000C3018614004200040607FE0844800000000001555155555FF";
    attribute INIT_27 of inst : label is "108008A100868002000020241020850045050000FFFFFFC00000000800C00C00";
    attribute INIT_28 of inst : label is "001980C4067831018CA90006218616B501111A550000000000E1C38304000028";
    attribute INIT_29 of inst : label is "002A00054002000150002A000540002800140001401500148052804A80295500";
    attribute INIT_2A of inst : label is "A801540002A0015400AA00015000AA00550000A80055002A800054002A801540";
    attribute INIT_2B of inst : label is "A0001550000A80001540002A8000540000AA001540000A80055002A800054002";
    attribute INIT_2C of inst : label is "B6893F91882F1551AD8C593B6B6FFE512EEF1BB3BFA69BB3BADBFF91FFD5000A";
    attribute INIT_2D of inst : label is "77608C1286736D6CDB92CE4B6E4D9BCE622763E430E318301906180EC7CCE1ED";
    attribute INIT_2E of inst : label is "A6DDB6B6DB6F440CE6EC32DBD8C2C9EDB6DB363DB6DB6CF9B6CF9B0150F54087";
    attribute INIT_2F of inst : label is "003D83B4DDC5B6E76C309D9B6CCEE9D6D06DB6CDB5B6C6CCC36666DB768B6D9B";
    attribute INIT_30 of inst : label is "3FE0000003FE001555C000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "AAD5555DFF55B6FAABBFFFBB6AB5577FF556D564A41001010010001101100000";
    attribute INIT_32 of inst : label is "1AAAAD555211AAAAD5552010000D5550015AAB555AAAD55AAB556AAD55AAB556";
    attribute INIT_33 of inst : label is "FFFFF808BFFFFFFBFC90DB6DB6DA07FFFF910002AAAA8000030000103FF83DB4";
    attribute INIT_34 of inst : label is "DB6A3FFFFD997FFFFFFC807FFE281AAAFFF5AAAFFF494E66666590666666489F";
    attribute INIT_35 of inst : label is "220054422315120409C44F60E152DD0208FB666C42A809B88484FFFFFE666641";
    attribute INIT_36 of inst : label is "F058CC2033EA0E371999556499A62304612021D31CF8720409CC913962A8CD11";
    attribute INIT_37 of inst : label is "244F8D1A05B830CB706C7331A623019B6CE41BB7C25646541E18D8C4C1B08916";
    attribute INIT_38 of inst : label is "80D920205007A633643648C1F20402810706201D1122244488D11B226548A915";
    attribute INIT_39 of inst : label is "81324069240620310124000120008CA03801923884C9027256EB0A9C52322714";
    attribute INIT_3A of inst : label is "C090F7BF863DE63F7F1E63F7E3CC44C9192ACEC6CECECEDA821B6E2C81388138";
    attribute INIT_3B of inst : label is "3F00F983F207E43E43C83FBDE61FDEF31F8F843F1E10FC7843F1E10A04C7E63F";
    attribute INIT_3C of inst : label is "35BD2B6E96D616B5B9AF2F863F93FFFF80000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0872068B413EFABC3AAF9FCADD010F6C9401820C088C3E1E5E3F9787F2F170FF";
    attribute INIT_3E of inst : label is "04068000000002B1375958AD6630AC8721BAB081A5106E4872126CCD243927CE";
    attribute INIT_3F of inst : label is "F9BD4C480C30B37CED49ECDB9005B166321BA861736134FF6221E3D351DA4390";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "07FF90F0600180681101150322E0104047BFC87FFF807C1043FCC1A1F9C1F1BA";
    attribute INIT_01 of inst : label is "8C8C002040000B82800FFE54244420C34D80D9DD384FB04D6E0DB0172234E380";
    attribute INIT_02 of inst : label is "FFFE6550A12A8A8842A884C7898020AA80D480C0111000000800214109801607";
    attribute INIT_03 of inst : label is "0000004020100805004092492492049240924924924012A0280C809F06C4881B";
    attribute INIT_04 of inst : label is "4040000000010000000000000002000000000002804020100800000000402100";
    attribute INIT_05 of inst : label is "8000000000000000008000000000004000000000000000000800200000000000";
    attribute INIT_06 of inst : label is "0000000020004040000000000080010000000000000020000000000000000000";
    attribute INIT_07 of inst : label is "9000000000000400000000012000000000001000100000000000000000000000";
    attribute INIT_08 of inst : label is "0210000000000000000000000000000010010000080000000000000000044000";
    attribute INIT_09 of inst : label is "0000000000020080100000004000840000000000000040100000000000000000";
    attribute INIT_0A of inst : label is "0000084040000000000000000001000000000000000000000000000001040000";
    attribute INIT_0B of inst : label is "0000000000000000102000000000001020480040000000020000400000000000";
    attribute INIT_0C of inst : label is "0000000000000000002000000200008000000000800000001000008002400000";
    attribute INIT_0D of inst : label is "1111425090A42D328E12BCE082E11C05131C4F81190000000000000000800000";
    attribute INIT_0E of inst : label is "79F02210000BE6CB0081004121A9A9DDA0898F81014D464F90D2907C12290101";
    attribute INIT_0F of inst : label is "7DB95561110C3AADCE915573B4028453E1022C001002AC82FB3C68CA3ECA395E";
    attribute INIT_10 of inst : label is "489122044682490405A842A480142140840A830C242C22838F0031088500FEDB";
    attribute INIT_11 of inst : label is "28584308524970861013843086106C44209044444849126880A4122044B06812";
    attribute INIT_12 of inst : label is "68C53290C48622C5113264C98248ACB3632E443841A1858824480C127B24625A";
    attribute INIT_13 of inst : label is "1B449116164DC4491653B176B888B0BB88C37710891A12E2242488B190184142";
    attribute INIT_14 of inst : label is "43925A186B9632412208488224199DB284924992C9A496492C92593B20489125";
    attribute INIT_15 of inst : label is "449B4953146CB32C24E4B7764C8022480AA05C245E7336C94501C00C4445924B";
    attribute INIT_16 of inst : label is "E6266776114207611483128850C14E0C9218960884900B024852235D0255B286";
    attribute INIT_17 of inst : label is "0E4804FD9372881204824594BBB59320304680223A4DCA201049111192C9D90E";
    attribute INIT_18 of inst : label is "C492441122124B3146180124A424922492329520529594844451B046493448E4";
    attribute INIT_19 of inst : label is "F60EC9D8848136A698242461020C49109225925CB54093180A301324901A0044";
    attribute INIT_1A of inst : label is "2493734926C60D90E4E404F240C960CAC250440C64B8B325F92E4C02CE4A226D";
    attribute INIT_1B of inst : label is "891D9C08433177F6DFDFE7209249249244832DF120010C126601200118040802";
    attribute INIT_1C of inst : label is "B484CC11DF77B2CB28089FF9AB12482421302C402010401A135588D111122E90";
    attribute INIT_1D of inst : label is "0028888ACED22220614610652404B68AB412B1F08960B580FFFFFE68F000000D";
    attribute INIT_1E of inst : label is "84444803C7081E38403C70818078E103041250504908B60C9106062888912224";
    attribute INIT_1F of inst : label is "A81025C4896D4200010898020444E1FE410424B648D1A068D034083A4F325927";
    attribute INIT_20 of inst : label is "2C99889105009408D21125B8000004F1EC2C16A58964920C48B24B2030946485";
    attribute INIT_21 of inst : label is "048C0C12C5227AFC849750B24CDEBB35B65B69B431CB52D2D1D0C888D2232CA2";
    attribute INIT_22 of inst : label is "1331213424889250D0D09BB1AF9883106F044998DF2419516C9A3692C918588A";
    attribute INIT_23 of inst : label is "85864332793180444207044042203444809B20D6E409F91B23686C4206724122";
    attribute INIT_24 of inst : label is "1010041000410040FFFFFFFB027F26A88D4262E071CC96C96D62C0C858642C0C";
    attribute INIT_25 of inst : label is "FE00000005555555504455557FFFFFFF7003800842000001090800420C000002";
    attribute INIT_26 of inst : label is "E11204895406006030C06154042AA0419FFF80844800000800001555555555FF";
    attribute INIT_27 of inst : label is "1000000102040000000000041000855000005000FFFFFFF80000C3B006006000";
    attribute INIT_28 of inst : label is "001928C3065230C196A94A18400008429422520000000000038706081C000000";
    attribute INIT_29 of inst : label is "00200004000200010000200004000020001000014A800014A900004A95000000";
    attribute INIT_2A of inst : label is "0001000002000100008000010000800040000080004000200000400020001000";
    attribute INIT_2B of inst : label is "0000100000080000100000200000400000800010000008000400020000040002";
    attribute INIT_2C of inst : label is "9288FF81902E05518DCE496B496FFF510DA619111F924B93BA5BF501FFC00008";
    attribute INIT_2D of inst : label is "F6208C0681512426D990EE43264993CE422E61C430A1183819071C0647CCE1E4";
    attribute INIT_2E of inst : label is "025D921249260248C26E3ACADCE2DDEC904B366D94D96648A6648A5400E04086";
    attribute INIT_2F of inst : label is "002DC1B459C492666E39D9DB26EEDD92502512CC9092424C8126425936012489";
    attribute INIT_30 of inst : label is "001FF0000001FF1555D555555555555555555555555555555555555500000000";
    attribute INIT_31 of inst : label is "AAD5D5555555B6DAAAAABAAB6AB555557556D574801110011100001110000000";
    attribute INIT_32 of inst : label is "35555AAAAA515555AAAAA515555AAAAA515AAB555AAAD55AAB556AAD55AAB556";
    attribute INIT_33 of inst : label is "00000C28C000000602946DB6DB6D4C2108430000000000008700001860043B6C";
    attribute INIT_34 of inst : label is "B6DA700003BBC00000029460000D3D550007D550006106EEEEEFB0EEEEEEDDB8";
    attribute INIT_35 of inst : label is "6A00D486A335220C010C5F60C3525C2410596E5806BA88904442FFFFFEEEEEC3";
    attribute INIT_36 of inst : label is "E0594C20032E04170B0955401084612C2500054218D0220C0104023962A0E035";
    attribute INIT_37 of inst : label is "00CD061C1DBC307B786C21108461228D6C440B6302D746D40C08C945C0A18B56";
    attribute INIT_38 of inst : label is "805000604006841125125848A20C0281450A203C300600C0184309602D01A034";
    attribute INIT_39 of inst : label is "802AC008A4002003002200000000880230010010008B0176D6AA1A8856B6A204";
    attribute INIT_3A of inst : label is "0000000002000000000020000004020401628AA08AA88ABA8209260D80298029";
    attribute INIT_3B of inst : label is "0000008001000200200400000200000100000000000000000000000000400000";
    attribute INIT_3C of inst : label is "38952B2696525294ACA7278617A0FFFF80000000000000000000000000000000";
    attribute INIT_3D of inst : label is "08522403001AA2AC2A0E9ED2491106949C05825C08DC3A1E4E179382F271227E";
    attribute INIT_3E of inst : label is "04008000000002B0A55950AC2220A40203AAA18087006440203064C40414068A";
    attribute INIT_3F of inst : label is "FC9B5C482491907CF64BC9C9900C91223249A823306102FF6200A1D351424290";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
