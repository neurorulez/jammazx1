-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0B92300C0C481F961DD41F96273C033012301F960B931DDD303835350F611A1C";
    attribute INIT_01 of inst : label is "AAAA000000005555444C000031110000000080CC000033020FC316340FC41796";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF0000000043C1182443C11824CC00CC0000330033";
    attribute INIT_03 of inst : label is "182482826559300C25582008241800007FFDB7FE7FFDB7FE7FFDB7FEFBEFC283";
    attribute INIT_04 of inst : label is "428118240960200824180000241800000960200842811824080C32061028B084";
    attribute INIT_05 of inst : label is "668918240AA00AA0C3C33EBCEC3B1694D0071694728D382C4FF1182442811824";
    attribute INIT_06 of inst : label is "123020081DD42A282BA92A280F78022031342A2813362AAA30302A2A0FC32028";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF1F9728281E9C2A28";
    attribute INIT_08 of inst : label is "0DD1222A1DD408801D1C2A2A0FC328A80CC022281FD62AA80FC30A8200000000";
    attribute INIT_09 of inst : label is "0FC32A283FDF0A823FFF0A820C0C2A2A3CE40AA203032A2830302A2A1FD70A82";
    attribute INIT_0A of inst : label is "3FD70A820FD720000FC32A28303020201D942A280FD30AA20FC3282A0FC30880";
    attribute INIT_0B of inst : label is "1004000000FF00FF00FF00FF00FF00FF00FF00FF32342AAA1B1E20203A3C0A82";
    attribute INIT_0C of inst : label is "0000100400FF00FF00FF00FF000000000000382C00FF00FF00FF00FF10040000";
    attribute INIT_0D of inst : label is "00FF00FF00FF00FF00FF00FF382C00000000000000FF00FF00FF00FF3EBC0000";
    attribute INIT_0E of inst : label is "4000000000FF00FF00FF00FF0000000044C0000000FF00FF00FF00FF00FF00FF";
    attribute INIT_0F of inst : label is "00FF00FF00FF00FF00FF00FF313400000000000000FF00FF00FF00FF33370220";
    attribute INIT_10 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_11 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_12 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_13 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_14 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_15 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_16 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_17 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_18 of inst : label is "13337FFFFFFFFFFF12E6CC009B840033884429991122666802FF00FF00000000";
    attribute INIT_19 of inst : label is "FCFCF3F37CFC0000FBFFFFFF0000C0C0000000003B3F0203FCECC080CCC4FFFD";
    attribute INIT_1A of inst : label is "00000000ABAB0000FBFFDFBFCFCFCCCC3F3FCFCFEAEA0000FFFBFCFFF3F33333";
    attribute INIT_1B of inst : label is "00FF00FF00FF00FF00FF00FF20DFF501112CF3F93D3F0000FBFFFFDF00000703";
    attribute INIT_1C of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF02FF00FF02FF00FF";
    attribute INIT_1D of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF08FF00FF08FF00FF";
    attribute INIT_1E of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF02FF00FF02FF00FF";
    attribute INIT_1F of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF08FF00FF08FF00FF";
    attribute INIT_20 of inst : label is "382CBBF54000000000008000C0C00000B554950F24B08643C52C20AFD643C12F";
    attribute INIT_21 of inst : label is "00000333331B00000000CCC0E4CC0000382CBBF543210000000080000C480000";
    attribute INIT_22 of inst : label is "01013BAF372C3333CFF0BFF738D8C0800323133320090000C8C0CCC460080000";
    attribute INIT_23 of inst : label is "2333FFFB15570323CCC0EFFFD554C8C001013BAD241C3333CFF08FDF3014C080";
    attribute INIT_24 of inst : label is "3031FFFB195F03234C0CEDFFF564C8C03031FFFB195F03234C0CEDFFF564C8C0";
    attribute INIT_25 of inst : label is "30303330000000000C0C0CCC000000000203333300000000C080CCCC00000000";
    attribute INIT_26 of inst : label is "0008313E031300002000BC4CC4C0000000303334010100000C001CCC40400000";
    attribute INIT_27 of inst : label is "03231BB33F7E0000C8C0CEE4BDFC00000323EDDF37350000C8C0F77B5CDC0000";
    attribute INIT_28 of inst : label is "0323133320090000C8C0CCC46008000003231333E8C90000C8C0CCC4632B0000";
    attribute INIT_29 of inst : label is "07029CDA09B82A952644D4FA95264494FA95264454FA9526641FF501112CF3F9";
    attribute INIT_2A of inst : label is "0D93CBF5CF08BCA3C0BBFAD0C7F72051FDD50954954955A5559087DE3B21FE0B";
    attribute INIT_2B of inst : label is "014000006A478D3491234504212375C421234504212E4504212E45042E4F1314";
    attribute INIT_2C of inst : label is "00000140421607DE421607DE0000000000000BE00EFFFF206451202901400000";
    attribute INIT_2D of inst : label is "5E7891235D6421141470860B0BE0000000000000134908481349F7902FF80000";
    attribute INIT_2E of inst : label is "400000002BAD8A245245659900000000740000009D49205245658959569A05A6";
    attribute INIT_2F of inst : label is "945D22D5D748B5A5D22C457701F400000000000015852099B046ECD401FF0028";
    attribute INIT_30 of inst : label is "6F411492B34DE152B34D2548B975522E69559B5B5566D45548A5155E6A49549A";
    attribute INIT_31 of inst : label is "415798D5515E6055CA05798557186558B5555E6E4974BB935D2ED4175AB5B5D2";
    attribute INIT_32 of inst : label is "0B34ACD21B8223B8A26B9A655981451566351CA056985471B15A6351C2395662";
    attribute INIT_33 of inst : label is "09616CB146E1E34D26C1B16EEC1BB359CEE22C18B34255E49669E496E9A69A69";
    attribute INIT_34 of inst : label is "556645942AC5A8863420AC13B6382A8A090860F095E65510A0AE2185E14822EC";
    attribute INIT_35 of inst : label is "14D27AEEFCB3428C1346082B04EE8E089082421B3C245599D0415E6559569958";
    attribute INIT_36 of inst : label is "B07BA4D1C13492090AC137956645104E288B06C5A69EB2C717DE47175C48A187";
    attribute INIT_37 of inst : label is "CB169DC2C135AD555999442C1060E68A411C13492191AC1379566551073C20B8";
    attribute INIT_38 of inst : label is "007F7FFFFFFFFFFF316ACC00A94C003399002A95006656A8A6D1369200000000";
    attribute INIT_39 of inst : label is "FFF0F0FF7FF00000FBFFFFFF0000F000000000000BFF000BFFE0E000FD00FFFD";
    attribute INIT_3A of inst : label is "00000000AAAF0000FBFFEF7FFF0FFF000FFFFF0FFAAA0000FEFFFFF3F0FF00FF";
    attribute INIT_3B of inst : label is "EF1AE21934EF4A749F72D64D5393C4C50364F2FD0FF70000FBFFFFDF0000040F";
    attribute INIT_3C of inst : label is "B4934EF4AB59354956702615CAE4E09853398573892B94DD27DD04B593549519";
    attribute INIT_3D of inst : label is "99F53333B7BA594DFFFCEFFFCA1B8E0B8A4E7C1C341CD749F766AE2EDA5EE51F";
    attribute INIT_3E of inst : label is "FFD46F410B07054CB12175C43AC485F79CB0623E2FEBFB272CB05F9764A51F64";
    attribute INIT_3F of inst : label is "800BC2FAE23C2FFFFCA7A0AD4D411818A0A4D08086068B06D508087510FF091B";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "1555302411142FE91554030311101FF5151523291514363C1010303010140FC3";
    attribute INIT_01 of inst : label is "AAAA00000000555540CC0000330100000000888C0000322215142B2B14143979";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF00000000241883C2241883C2CC00CC0000330033";
    attribute INIT_03 of inst : label is "41412418300C9AA610041AA4000018243D7CFFBF3D7CFFBF3D7CFFBF3D7CE3CB";
    attribute INIT_04 of inst : label is "241881421004069000001824000018241004069024188142604C3010210D1408";
    attribute INIT_05 of inst : label is "24189946055005503D7CC3C32968DC372968E00B341CB14E24188FF224188142";
    attribute INIT_06 of inst : label is "2FEB300C262C0FC32EE8074333342BBA2B3A07432F692C6C3034303025380F86";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF2F6903122D6823E3";
    attribute INIT_08 of inst : label is "262E0F872EEA0CC02E2E0C0C2DF80FD2272D0D852FE90FC3253C2FEB00000000";
    attribute INIT_09 of inst : label is "2F690FC30FC72FF30FD72FC30C0C0C0C0FD23DF8030307433A3A30300FC30FC3";
    attribute INIT_0A of inst : label is "0FC32FFF0FC33A3C0FC30FC33A3A30302D7807432FE93DF82F692FF22FE92EE8";
    attribute INIT_0B of inst : label is "0000200800FF00FF00FF00FF00FF00FF00FF00FF2BBB2C4C0F0F30300FD72F7D";
    attribute INIT_0C of inst : label is "0000000000FF00FF00FF00FF000000000000100400FF00FF00FF00FF00002008";
    attribute INIT_0D of inst : label is "00FF00FF00FF00FF00FF00FF100400000000000000FF00FF00FF00FF3D7C2008";
    attribute INIT_0E of inst : label is "0000800000FF00FF00FF00FF00000000000088C000FF00FF00FF00FF00FF00FF";
    attribute INIT_0F of inst : label is "00FF00FF00FF00FF00FF00FF000032380000000000FF00FF00FF00FF0110333B";
    attribute INIT_10 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_11 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_12 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00DD00FF00FF00FF00DD00DF";
    attribute INIT_13 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_14 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_15 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_16 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_17 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_18 of inst : label is "0103373FFFFFFFFF1666448899942211CC0021D90033674800FF00FF00000000";
    attribute INIT_19 of inst : label is "CCCCF3F3CFFF8888BCFCFFEF0000000000000000BFFF2333FFFECCC8C040FCDC";
    attribute INIT_1A of inst : label is "00000000FFEF0202C0C0FDFFCFCFCCCC3333CFCFF3FF80800303FFF7F3F33333";
    attribute INIT_1B of inst : label is "00FF00FF00FF00FF00FF00FF30E386E42A44FD11FFF722223F2FF3EF00000000";
    attribute INIT_1C of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_1D of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_1E of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_1F of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_20 of inst : label is "0CB0D4D0022200000000C0C0C8C00000BFD050CB08D0DE32C634378469F2C21E";
    attribute INIT_21 of inst : label is "0203333300010000C080CCCC782C00000FB0D4D2213800000000C0C00C8C0000";
    attribute INIT_22 of inst : label is "03207FF400002303E1735CED0000CCC03033031300000000CC0CC4C0382C0000";
    attribute INIT_23 of inst : label is "2BBFFBFF00003333FEE0FFCF0000CCCC032077FD00002303E1730E790000CCC0";
    attribute INIT_24 of inst : label is "389CFD3F00003033362CFAFF0000CC0C389CFD3F00003033362CFAFF0000CC0C";
    attribute INIT_25 of inst : label is "323C0313000000003C8CC4C0000000002333031300000000CCC8C4C000000000";
    attribute INIT_26 of inst : label is "320F333400000000F08C1CCC00000000303C1313000000003C0CC4C400000000";
    attribute INIT_27 of inst : label is "30337DEF11100000CC0CFB7D0444000088F33EFC00000000CF223FBC00000000";
    attribute INIT_28 of inst : label is "30330313382C0000CC0CC4C0382C0000303303137F7E0000CC0CC4C0BDFD0000";
    attribute INIT_29 of inst : label is "020201D308E634955398C644955398C644955398C6449553B8E386E42A44FD11";
    attribute INIT_2A of inst : label is "44013154840AE6F1069E5F4EA864742BCC0F0874E75F9DBE74F3C3CCBFAA190B";
    attribute INIT_2B of inst : label is "0000028029AFC4412B3100082B3118682B3108282B3310482B370008212456AA";
    attribute INIT_2C of inst : label is "0000000082B3118682B7110400000000000001409ACCCCB9A66AB9AD00000280";
    attribute INIT_2D of inst : label is "9248EB3310482B004788DA1B014000000000000044120ACCC00254871FF40280";
    attribute INIT_2E of inst : label is "00008000959649219E79E78A000000000000B8009A59E19249A48A79E59E2924";
    attribute INIT_2F of inst : label is "60115769C455DA6111369444000002F80000000074DD30994582F120001402FF";
    attribute INIT_30 of inst : label is "769074C0C49D7340C49D7555D631557588545DA31517680544DA11513584544D";
    attribute INIT_31 of inst : label is "84554EA011553B80638554E6018DA555DA01513780454DE41153790455DE5115";
    attribute INIT_32 of inst : label is "2C49ADD779DE76ADAF79CE3554EE311553B8C638554EA318E155388C63695138";
    attribute INIT_33 of inst : label is "9D2D264582FBF11049164591116CC49961109166C48255E792792696ED869969";
    attribute INIT_34 of inst : label is "1513684A731530DA05E6B166B169A1E3698DAEC0951378863680369D374C2111";
    attribute INIT_35 of inst : label is "11C7B130C2C48220D05E79AC59AC5A6979DA636AB024544D2011513788544D20";
    attribute INIT_36 of inst : label is "C58CA41BC010637B7B1674D553780742302C591696D38EEF10C3AF10C38DE7AF";
    attribute INIT_37 of inst : label is "245A913B1674D16544DE00B1674023884DBC000237B7B1674D55368077B16AC6";
    attribute INIT_38 of inst : label is "000707FFFFFFFFFF156A6600A9540099CC0032950033568CB51E74D300000000";
    attribute INIT_39 of inst : label is "FF00F0FFFF3FAA00BFF0FFEF0000000000000000BFFF00BFFFFEFE00D000FFD0";
    attribute INIT_3A of inst : label is "00000000FFEF000AF000FFF7FF0FFF0000FFFF0FF3FFA000000FFDFFF0FF00FF";
    attribute INIT_3B of inst : label is "5C49034875A35A7DB2CCF2CB34E3B5281988CCD5FDFF00AA0FEFF3EF00000000";
    attribute INIT_3C of inst : label is "58D75A35A3CB2CD2C76075D71A35A1D75C0D75C69D68D71F6CB82B3CB2CD2C15";
    attribute INIT_3D of inst : label is "46F4888835D14D157331A7331A49DA49DA88FC8B20A807DB2C199D512749959C";
    attribute INIT_3E of inst : label is "A95DE21A6C5A1A43BB310C380EECC430E2C5A0BD3BDAF678B0458CF14C402FCC";
    attribute INIT_3F of inst : label is "2A5B165F0AB1673332FCE1E21A0D7B79EDE017B79EDE2C59167B78059FCC1E6A";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "1FD7300C191C0FC31DD40B833338177517350B831F961C9C303830301A340F49";
    attribute INIT_01 of inst : label is "AAAA000000005555404C0000310100000000808C000032021F9603211E9413D3";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF00000000000000000000000000000000CC00CC0000330033";
    attribute INIT_03 of inst : label is "012DB4800000000000000000000000003FFCD3B33FFCD3B33FFCD3B3BFFE7FFD";
    attribute INIT_04 of inst : label is "0000000000000000000000000000000020081004382C341C49618692484C3212";
    attribute INIT_05 of inst : label is "269819640FF00FF03EBC3D7C3EBC3D7C3EBC3D7C382C341C382C341C382C341C";
    attribute INIT_06 of inst : label is "0761300C0C842F692EE82F691B3C033021302F6907632EEE30343A3A0F92252C";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF0FC329380FC82B69";
    attribute INIT_08 of inst : label is "0C84272F0CC00CC00C0C2E2E0FD22DF80D85272D0FC32FE90F960FC300000000";
    attribute INIT_09 of inst : label is "0FC32F692FCF0FD32FFF0FC30C0C2E2E2DF01FF203032F6930303A3A0FC30FC3";
    attribute INIT_0A of inst : label is "2FC30FD70FC330140FC32F69303030300DD02F690FC31FF20FC32D7A0FC30CC0";
    attribute INIT_0B of inst : label is "0000000000FF00FF00FF00FF00FF00FF00FF00FF23312EEE0F0F30302F7D0FD7";
    attribute INIT_0C of inst : label is "0000000000FF00FF00FF00FF000000000000382C00FF00DD00DD00FD00000000";
    attribute INIT_0D of inst : label is "00FF00FF00FF00FF00FF00FF382C00000000000000FF00FF00FF00FF3FFC0000";
    attribute INIT_0E of inst : label is "0000000000FF00FF00FF00FF000000000080004000FF00FF00FF00FF00FF00FF";
    attribute INIT_0F of inst : label is "00FF00FF00FF00FF00FF00FF202010100000000000FF00FF00FF00FF23321331";
    attribute INIT_10 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_11 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_12 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_13 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_14 of inst : label is "00FF00FF00FF00FF00FF00DF00FF00FF00FF00DD00DD00DD00DD00FD00FD00FD";
    attribute INIT_15 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_16 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_17 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_18 of inst : label is "03233FBFFFFFFFFF16E6CC009B940033CC0029D90033676800FF00FF00000000";
    attribute INIT_19 of inst : label is "ECECF3F3000080800000000000000000000000003F7F0313FDFCC4C0C8C0FEFC";
    attribute INIT_1A of inst : label is "000000000000ECEC15150000CFCF7F7F3B3BCFCF00003B3B54540000F3F3FDFD";
    attribute INIT_1B of inst : label is "00FF00FF00FF00FF00FF00FF12D5666695555955000002020000000000000000";
    attribute INIT_1C of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FD00DD00DD00DD00DD00FD00DD00FF";
    attribute INIT_1D of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_1E of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_1F of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_20 of inst : label is "0102CCC00000373EFFDCFEDBE0E0D8CC633EAAD103C8EBB64CF23AC095B45089";
    attribute INIT_21 of inst : label is "7BDEE4CC28081233BFFD323B302CCCC40002CCC00330373EFFDCFEDB2C2CD8CC";
    attribute INIT_22 of inst : label is "363E000000032323C8C00000C000C4C04CCCF7DF220A13313331F7EFB08CCC84";
    attribute INIT_23 of inst : label is "0001033320221332400CCCC08C0C8CC4363E000003302323C8C070000C0CC4C0";
    attribute INIT_24 of inst : label is "2333000030301233CCC800000C0CCC842333000020201233CCC800000C0CCC84";
    attribute INIT_25 of inst : label is "3337233300000001DCCCCCC8000040000313233300000000C4C0CCC800000000";
    attribute INIT_26 of inst : label is "323E333F02021332BC8CFCCC8080CCC41335333300003137DCC4CCCC0000DC8C";
    attribute INIT_27 of inst : label is "4CCCFFDF3B3A13313331F7FFACECCC8434CCBFFF22203137233CFFFE0888D8CC";
    attribute INIT_28 of inst : label is "4CCCF7DF320E13313331F7EFB08CCC844CCCFFDFFFFF03333331F7FFFFFFCCC0";
    attribute INIT_29 of inst : label is "43D131E344F83BD203309AEBD203309A6BD203309AABD2031295666695555955";
    attribute INIT_2A of inst : label is "62762602E2AD353AA2E363E4DEC130064C50461AC18C063019CB2B64BD379046";
    attribute INIT_2B of inst : label is "01400000C11B48964613114116122591161211411613218116130101128A85F4";
    attribute INIT_2C of inst : label is "0000014011693010116130100000000000000BE0E9EEEE4E848C4E9D01400000";
    attribute INIT_2D of inst : label is "20B3C613218116209C20E3260BE0000000000000C0404584C040985B2FF80000";
    attribute INIT_2E of inst : label is "40000000082482CF28B20B38000000007400000028928D2092C930824B24D28B";
    attribute INIT_2F of inst : label is "825E03305780CC05ECB3097A01F40000000000007ADA345E2B118AC801FF0028";
    attribute INIT_30 of inst : label is "710168E0AB1E36A0AB1E3480F415203D014A0F815283E014B2F825283F0D490F";
    attribute INIT_31 of inst : label is "0D4A0C436D28300D8334A0C4360E34A2FC25243C017B0C435EC310D782C405EC";
    attribute INIT_32 of inst : label is "0AB299E3A4E93A7E9F04C1F480C836D20300D833480C0360DD20330D83AD2C30";
    attribute INIT_33 of inst : label is "1E1E386B11F6D22590AC6B39AACA2B1E02AC2AC8AB114AD869A65B6D8A38A182";
    attribute INIT_34 of inst : label is "5243F099391A98E31A9ACAC8418E11338D8E34A4D283E05938EE38DE368D1398";
    attribute INIT_35 of inst : label is "029A281A806B118021A9A6B2B21063844CE3638D19334B0F815D283E05480F81";
    attribute INIT_36 of inst : label is "2B243866481443A7AEAC78D283C055913F22B2AC0821419900511900100E5959";
    attribute INIT_37 of inst : label is "6AB0AB1AAC78CAC490FC160AC58D1370826480403A7AEAC78D283D05593AFEA4";
    attribute INIT_38 of inst : label is "007F7FFFFFFFFFFF316ACC00A94C003399002A95006656A828A078CD00000000";
    attribute INIT_39 of inst : label is "FFF0F0FF0000F0000000000000000000000000000BFF000BFFE0E000FD00FFFD";
    attribute INIT_3A of inst : label is "000000005500FFF000000000FF0F0FFF0FFFFF0F00550FFF00000000F0FFFFF0";
    attribute INIT_3B of inst : label is "829EE39E1E31E31C71DC71C7B80801FF901509000000000F0000000000000000";
    attribute INIT_3C of inst : label is "A0F1E31E31C71EE4C3EC3E29213E14F8A80F8A484F84F8071C7B031C71EE4C03";
    attribute INIT_3D of inst : label is "48D6EEEE1E00CF9AFBBA37BBA39423942339B41AEC07E1C71DA6A2EEE3D93522";
    attribute INIT_3E of inst : label is "02667364EAB3E43066100103C598401446AB1CD2312C43A0AA2B28BB58744DD8";
    attribute INIT_3F of inst : label is "72B5AF23DC9AF3BBB934CE726482A7AE5E786A7AE5E76AB0AC979D792F224DAA";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0110302404403FBC1554171605140BB01010373C0111377D1010353505411A96";
    attribute INIT_01 of inst : label is "AAAA00000000555544CC000033110000000088CC0000332205413E3E05443D3C";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF00000000000000001004200800000000CC00CC0000330033";
    attribute INIT_03 of inst : label is "3008100C1004200810042008100420087D3DAF7A7D3DAF7A7D3DAF7A796DB7DE";
    attribute INIT_04 of inst : label is "000000000000000000000000100420081414282815542AA810042008200C3004";
    attribute INIT_05 of inst : label is "640998060000000015542AA815542AA815542AA815542AA815542AA815542AA8";
    attribute INIT_06 of inst : label is "3ABA2008377C0A822BA9020227702AAA3B3E02023B3C28283030202025690A82";
    attribute INIT_07 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF3F3D02023C3C22A2";
    attribute INIT_08 of inst : label is "277B0A823FFE08803F3E08082DE90A82266808803FFC0A8225692AAA00000000";
    attribute INIT_09 of inst : label is "2F690A821FD72AA21FD72A820C0C08081EC628A8030302023A3A20201FD70A82";
    attribute INIT_0A of inst : label is "1FD72AAA0FD72A280FC30A823A3A20203D3C02022FF928A82F692AA22FE92AA8";
    attribute INIT_0B of inst : label is "1004200800FF00FF00FF00FF00FF00FF00FF00FF3ABE28081B1E20201A962A28";
    attribute INIT_0C of inst : label is "0000100400FF00FF00FF00FF000000000000100400FF00FF00FF00FF10042008";
    attribute INIT_0D of inst : label is "00FF00FF80FF00FF00FF00FF100400000000000000FF00FF00FF00FF3C3C2008";
    attribute INIT_0E of inst : label is "4000800001FF11FF00FF00FF000000004440888010FF00FF00FF00FF01FF10FF";
    attribute INIT_0F of inst : label is "00FF00FF00FF00FF00FF00FF111422280000000000FF00FF00FF00FF1115222A";
    attribute INIT_10 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_11 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_12 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_13 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_14 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_15 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_16 of inst : label is "00FF00FF11FF10FF00FF00FF01FF01FF00FF00FF11FF00FF00FF00FF00FF10FF";
    attribute INIT_17 of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_18 of inst : label is "1113777FFFFFFFFF1266448899842211884421991122664800FF00FF00000000";
    attribute INIT_19 of inst : label is "DCDCF3F300004040000000000000000000000000BBBF2223FEEEC888C444FDDD";
    attribute INIT_1A of inst : label is "000000004444DCDC2A2A0000CFCFBFBF3737CFCF11113737A8A80000F3F3FEFE";
    attribute INIT_1B of inst : label is "00FF00FF00FF00FF00FF00FF00C0111501510004000001010000000000000000";
    attribute INIT_1C of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_1D of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_1E of inst : label is "00FF00FF01FF10FF00FF00FF01FF00FF00FF00FF00FF11FF00FF00FF00FF01FF";
    attribute INIT_1F of inst : label is "00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF";
    attribute INIT_20 of inst : label is "020180C04222233BEEB4CFFDDDC4E8E02FFC4FC1401CDCF05007370F71F0500B";
    attribute INIT_21 of inst : label is "B9BDDCCC0444232B5E6E33373938E848000180C26129233BEEB4CFFD1DCCE8E0";
    attribute INIT_22 of inst : label is "0981444202233313C4408100C080C880988C6FE71515032B3026FBF97C7CE8C8";
    attribute INIT_23 of inst : label is "00122323111123218400C8C86CCC48C80981444221293313C44080800CC8C880";
    attribute INIT_24 of inst : label is "1033000022282123CC8400002888C8481033000000002123CC0400002888C848";
    attribute INIT_25 of inst : label is "333B131300000202ACCCC4C4000080802223131300000000C888C4C400000000";
    attribute INIT_26 of inst : label is "312D32360111222A784C9C8C4440A888233B131701012333ECC8D4C44040CCC8";
    attribute INIT_27 of inst : label is "988C6FEF1555232B3026FBF95554E8C8BC8C7FFF15152B3B323EFFFD5454ECE8";
    attribute INIT_28 of inst : label is "988C6FE73D3D032B3026FBF97C7CE8C8988C6FEF7F7F232B3226FBF9FDFDE8C8";
    attribute INIT_29 of inst : label is "031C3CF04030340B0021C0740B0021C0740B0021C0740B0000C0111501510004";
    attribute INIT_2A of inst : label is "555545574F3BD7D3C08D4D7C6441E03B4C3F730E30D3C30F0C33CC303F191272";
    attribute INIT_2B of inst : label is "00000280C32F04514B001451CB001C71CB001451CB031041CB431041C5455400";
    attribute INIT_2C of inst : label is "000000001CB001C71CB001C700000000000001405C333335C1C835C400000280";
    attribute INIT_2D of inst : label is "14500B031451CB010200DC420140000000000000041072D004103DC71FF40280";
    attribute INIT_2E of inst : label is "00008000041041021C71C704000000000000B800186183186146085145141145";
    attribute INIT_2F of inst : label is "840B002102C00850B002182C000002F8000000002C0B470BB710ADC3001402FF";
    attribute INIT_30 of inst : label is "02142D0F770F00CF770F02C00840B002142C00450B001182C00860B002182C00";
    attribute INIT_31 of inst : label is "182C004400B001100302C004400DC2C00850B0021C2C00850B002142C00860B0";
    attribute INIT_32 of inst : label is "477188F06018460184501402C008500B002140302C008500C0B002140370B002";
    attribute INIT_33 of inst : label is "0D41407710CBC11453DCB72EEDCBF70B2EF01DC0771C3DC71C6185148B2CB2CB";
    attribute INIT_34 of inst : label is "0B00210033CF3CDC0DC73DC70371C343700DC4750B002144370B370B02D1C3FC";
    attribute INIT_35 of inst : label is "01C720EC30771C1C30DC71CB71C0DC70C0DC03701D482C00C620B002142C00C4";
    attribute INIT_36 of inst : label is "770F2C3B4041047073DC3C0B003143D0000773DC3CB71CAD01C72D01C711C72D";
    attribute INIT_37 of inst : label is "0770B1E1DC3C3D42C00C421DC3F10003C3B4041047072DC3C0B003143C1DC87C";
    attribute INIT_38 of inst : label is "000707FFFFFFFFFF156A6600A9540099CC0032950033568C2FDC3C0300000000";
    attribute INIT_39 of inst : label is "FF00F0FF00000000000000000000000000000000BFFF00BFFFFEFE00D000FFD0";
    attribute INIT_3A of inst : label is "000000000000FF000FFF0000FF0FFFFF00FFFF0F000000FFFFF00000F0FFFFFF";
    attribute INIT_3B of inst : label is "335073531D81D81C71C071C73551550015555155000000000000000000000000";
    attribute INIT_3C of inst : label is "2071D81D81C71CD4F1F21CF2D81D8873CB873CB6076073C71C7C001C71CD4F87";
    attribute INIT_3D of inst : label is "000F33331CD2C7CB4CCD84CCD850D850D8CDC00F300C31C71CC88888B1FD1C73";
    attribute INIT_3E of inst : label is "00FDC71C47721C072B401C701CAD0071C0770012012449711F7734DD5C1C005C";
    attribute INIT_3F of inst : label is "1071DC4D041DC4CCCFDC21C71CC37071C1CC37071C1C0773D470731C7033CF73";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
