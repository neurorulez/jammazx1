-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "5555000003D5000057C00000015503C0554003C057D503C03C0F05783D0C255E";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF0000000033333333333333333333333303C003C0";
    attribute INIT_03 of inst : label is "3333333333333333333333333333333333333333C68325582828282807D027D8";
    attribute INIT_04 of inst : label is "3333333333333333333333333333333333333333333333333333333333333333";
    attribute INIT_05 of inst : label is "3333333333333333333333333333333333333333333333333333333333333333";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333332D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "FFFF2FF81E3450448D1410848DD710848D14108401F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "8940000857D70000460810900018014057D503C07FFD03C0FFFF2FF8FFFF2FF8";
    attribute INIT_0D of inst : label is "BD7E0000569503C0582503C0A00A0C3060090280182400000690000001602400";
    attribute INIT_0E of inst : label is "8142955621480AA01BE4000003C00D700C300960C003255807D0E00B55550000";
    attribute INIT_0F of inst : label is "1FF4028007D00000C0039556300C25580C300960055294009414001650050960";
    attribute INIT_10 of inst : label is "03C00BE00FF00000214828280820D007F82F3FFCE00BBD7E8002B41E7FFD0BE0";
    attribute INIT_11 of inst : label is "FFFFFFFF0000000000000000FFE0E000FD00FFFD00000000A940003E016ABC00";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000BFF000B007F7FFF";
    attribute INIT_13 of inst : label is "000AA00000000000000000000000000000000000000000000000000000000000";
    attribute INIT_14 of inst : label is "AAAA0000003C000000003C000000003C3C000000A000000A0A0000A000A00A00";
    attribute INIT_15 of inst : label is "34704D248A4AB255E7598545938A22C9B345052E49334C50364F39EF09600000";
    attribute INIT_16 of inst : label is "9D462B259839B1549A79604704D248E4EB255E75999459CF282E2C9ED549278E";
    attribute INIT_17 of inst : label is "E19BC4B261772C986F2C9B42F4A052CB75569209A0AD9BCB36D8F2C955AD1759";
    attribute INIT_18 of inst : label is "991459823B2C9820BB4514922861278EE820EED545268A1869E5BA08592C9B36";
    attribute INIT_19 of inst : label is "447B99F0493333B7BA59505C6ED1ED1DD5E749950598B2508AEC26DEC5455A75";
    attribute INIT_1A of inst : label is "541708EC22AA691890B989B7487B99F44967C1D41729F4E5F4E5342534255555";
    attribute INIT_1B of inst : label is "41519EF3A6239346F42749F72D64D505519F2A08AA4624239A62D0694BA51E17";
    attribute INIT_1C of inst : label is "EE59F949346F42B59354156702697C2E4609A5B39A5F1890B96DD27DD04B5935";
    attribute INIT_1D of inst : label is "6567FE5793333B7BA5945FFFC6FFFC23B862B824E7C1C341CD749F76E26A65A5";
    attribute INIT_1E of inst : label is "B2623E2FEBFB072CB25F9764A51F6499F5554575656565150525C5F5E59585B5";
    attribute INIT_1F of inst : label is "A4D28286068B26D108084590FF093BFCD46F490B270D4CB12175C43AC485F79C";
    attribute INIT_20 of inst : label is "3403E00307830082C01CC00BC2D0FA0012301F960B931DDD303835350F611A1C";
    attribute INIT_21 of inst : label is "B5001555017A000200545557AD4080000DF80C01017A02AA00E0F81C81F00000";
    attribute INIT_22 of inst : label is "00600C00005A000000C06030A400000002C30E83001F0000C780C2B041000000";
    attribute INIT_23 of inst : label is "00B3038300050000DE00C2C00400000003D00155001E000005C055F0B4000000";
    attribute INIT_24 of inst : label is "00B40055000500001E8057C050000000003500E0000000007800610000000000";
    attribute INIT_25 of inst : label is "002500C0000000005800610000000000003200E300000000F800CB0000000000";
    attribute INIT_26 of inst : label is "0020003300000000A000CC000000000000290015000000006800570000000000";
    attribute INIT_27 of inst : label is "002A000500000000A0005C0000000000002A0018000000008000610000000000";
    attribute INIT_28 of inst : label is "37F70CCC015F0000F7F7CCF3FD5000003FFFFFFF07FF00AFFFFCFFFFFFD0FA00";
    attribute INIT_29 of inst : label is "DFDF3333057F0000DF7F322BFD500000DFDF3333057F0000DFD733F9FD500000";
    attribute INIT_2A of inst : label is "0B4F08D000AF000BF1E00720FA00E000DFDF3333057F0000DFD7333CFD500000";
    attribute INIT_2B of inst : label is "002F08D007AF0002F8000720FAD080002C17FFD000080000E1E03FFD0D000000";
    attribute INIT_2C of inst : label is "98040200755F000E49334C50364F39EF9C17DFD007880000E8003FD400000000";
    attribute INIT_2D of inst : label is "9FF600006559300C4961300C82820C3042812008096000002418000010240480";
    attribute INIT_2E of inst : label is "9006955612842828396C0000300C1C340C301824C0031694341CC28355550000";
    attribute INIT_2F of inst : label is "3D7C2008341C0000C003955603C016940C301824141684408550011241411824";
    attribute INIT_30 of inst : label is "300C382C3C3C000012840AA00820C143CBE33FFCC2839FF6800287D27FFD382C";
    attribute INIT_31 of inst : label is "FFFFFFFF0000000000000000FCECC080CCC4FFFD000000009884033212268CC0";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000003B3F020313337FFF";
    attribute INIT_33 of inst : label is "0202808000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "AAAA00000330000000000CC0000003300CC00000808002020808202020200808";
    attribute INIT_35 of inst : label is "14F04D249A0A91D9D69D9505A24E328991CD072648375C1017CB3BE718240000";
    attribute INIT_36 of inst : label is "9D4609AD8A7191D49A79518334127920C9AD5D79A9547B470BA22F92D645278E";
    attribute INIT_37 of inst : label is "E297E43251B72E904FAC984EE4E0724B55D68249A3A1BA4F36D8F2C96765165D";
    attribute INIT_38 of inst : label is "895468460BEC886099CD245218A1278EC8A0FD9945268A1879A58AC84B64897E";
    attribute INIT_39 of inst : label is "5633B874483721FF9AD953507C99CF95F5676915261490D8BB28379AD5055979";
    attribute INIT_3A of inst : label is "45533B2022AA4A94A271A9375A33B9745927F114066DF5E1F5E105E105E15555";
    attribute INIT_3B of inst : label is "5015BC7B84AB914EC5E379371DA4C54563570A88998A04A3986AD261692D0D5B";
    attribute INIT_3C of inst : label is "DE99DAC517E36139915C156712294FE24609A4B79B5B28509BE5D379D2434975";
    attribute INIT_3D of inst : label is "55A7DDDB807F1AFFA5947F7FF73BCCE398E289E0F48DD00DDD349D7ED2AA65A5";
    attribute INIT_3E of inst : label is "90EA0FEBFABF072C93DB956C87976691D5D5553555A545950525F535E595A535";
    attribute INIT_3F of inst : label is "B492A10A260B34990A006414CECD3BFCD7634A07078D6C3111B5C632E501E7DC";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "0000000003C0000003C00000000003C0000003C003C003C005540AAF05501AF5";
    attribute INIT_02 of inst : label is "FFFFFFFF00000000FFFFFFFF0000000033333333333333333333333303C003C0";
    attribute INIT_03 of inst : label is "33333333333333333333333333333333333333331AA4C9431414141401401AA4";
    attribute INIT_04 of inst : label is "3333333333333333333333333333333333333333333333333333333333333333";
    attribute INIT_05 of inst : label is "3333333333333333333333333333333333333333333333333333333333333333";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333331EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "1FF4FFFFBF1145ACC40020ACC461A0ACC420A0AC2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "1000029100008280182004841AA403C003C003C007D02FF81FF4FFFF1FF4FFFF";
    attribute INIT_0D of inst : label is "D0070BE003C0A96A03C0A41A0C30500506902418014009600000028000240680";
    attribute INIT_0E of inst : label is "6AA9428105501284000027D80EB003C006900C301AA4C00300007EBD0000AAAA";
    attribute INIT_0F of inst : label is "01402FF800000BE06AA9C0031AA4300C06900C3000294AA0680028290690A00A";
    attribute INIT_10 of inst : label is "07D003C000000FF014141284E00B04107FFDF41F7EBDD007782D400107D0BFFE";
    attribute INIT_11 of inst : label is "FFFFFFFF0000000000000000FFFEFE00D000FFD0000000007C000295003D5680";
    attribute INIT_12 of inst : label is "0000FFFF00FF000000FFFFFF0000FF00FFFFFFFF000000FFBFFF00BF000707FF";
    attribute INIT_13 of inst : label is "000550000000000000FF00FFFF000000FFFF00FFFF00FFFFFF00FF00FFFF0000";
    attribute INIT_14 of inst : label is "0000555500003C00003C00003C0000000000003C500000050500005000500500";
    attribute INIT_15 of inst : label is "06F00418DEDEC5913554CE01508C0B1645A1B56380485281988CCC8D00000690";
    attribute INIT_16 of inst : label is "C6008C595C08E2159249236F00008DEDEC5913554C20152C5BB0B1602159249E";
    attribute INIT_17 of inst : label is "2214C245958591655191654245E08A9CC544D38D2091242459D23B1644D1A544";
    attribute INIT_18 of inst : label is "4CA015637BB16E3680865592323D249E327DE02195648C8F49248C9F4AB16459";
    attribute INIT_19 of inst : label is "44A659C78D888835D14D109920210211113554CA2152C5B8DE31A17316251354";
    attribute INIT_1A of inst : label is "31618D2634875959D58D476445A659C58DCFD084265834343434747474746444";
    attribute INIT_1B of inst : label is "D6C155C4903487563567DB2CCF2CB35B315C4A8D26567560D450829D8074BF10";
    attribute INIT_1C of inst : label is "9959C58D7563563CB2CD6C7607516163561D4580D45859D58D41F6CB82B3CB2C";
    attribute INIT_1D of inst : label is "866731E48888835D14D19733167331649D649D688FC8B20A807DB2C1D9511274";
    attribute INIT_1E of inst : label is "C5A0BD3BDAF668B0458CF14C402FCC46F4C4C4D4D4C4F4F4D4F4A494B494B4A4";
    attribute INIT_1F of inst : label is "A017B79ADA2C591A6B68259FCC1E6AA81DA21A6C5A1A43BB310C380EECC430E2";
    attribute INIT_20 of inst : label is "D0033803005F0B43C007C02C4100C1E0151523291514363C1010303010140FC3";
    attribute INIT_21 of inst : label is "EAAA6A00000102B5AAA800AD40005E80341F070000000F8180301F8055405E80";
    attribute INIT_22 of inst : label is "0C060300000000250030060000005A000D4301E300000082C170C3400000F800";
    attribute INIT_23 of inst : label is "0343007B00000020C1C0CD000000A0000FAA03A00000002DAA000BC000007800";
    attribute INIT_24 of inst : label is "03AA01780000000AAA002D000000A0000086001E000000000700AE0000000000";
    attribute INIT_25 of inst : label is "0086001A000000000300A4000000000000D3001F00000000C7004C0000000000";
    attribute INIT_26 of inst : label is "0033000500000000CC0004000000000000EA001600000000A800940000000000";
    attribute INIT_27 of inst : label is "003A000500000000A00054000000000000860001000000001800540000000000";
    attribute INIT_28 of inst : label is "0CCC3BFB000002AFCCF2FBEA0000FEA0FFFF3FFF005F0BFFFFFFFFFCF500FFE0";
    attribute INIT_29 of inst : label is "3333EFEF00000ABF3327EFBF0000FEA03333EFEF00000ABF339EEFAA0000FEA0";
    attribute INIT_2A of inst : label is "00B5004B001F00BF5E00E100F400FE003333EFEF00000ABF3396EFEB0000FEA0";
    attribute INIT_2B of inst : label is "00B5084B006B000B5E00E120E900E000FFE01C2B000000043FFED2D000000E00";
    attribute INIT_2C of inst : label is "004020190000A00380485281988CCC8DEFE06C2B00000B443FE8D40000000000";
    attribute INIT_2D of inst : label is "C143382C300C9AA6300C86920C30414124180690100418240000200801202408";
    attribute INIT_2E of inst : label is "6AA96009141421480000369C2C38300C24180C302968C00300006FF90000AAAA";
    attribute INIT_2F of inst : label is "10043EBC0000382C6AA9C003296803C024180C300221682848800AA124188282";
    attribute INIT_30 of inst : label is "341C300C00003C3C05502148C28304107FFDC7D36FF9C1434BE14001341CBFFE";
    attribute INIT_31 of inst : label is "FFFFFFFF0000000000000000FFFECCC8C040FCDC000000004CC0211903316448";
    attribute INIT_32 of inst : label is "0000FFFF333300003333FFFF0000CCCCFFFFFFFF00003333BFFF23330103373F";
    attribute INIT_33 of inst : label is "010140400000000033333333CCCC0000FFFF3333CCCCFFFFCCCCCCCCFFFF0000";
    attribute INIT_34 of inst : label is "0000555500000CC0033000000CC0000000000330404001010404101010100404";
    attribute INIT_35 of inst : label is "34380610FF5AE41515D4CC096340091E642594E792006049AB40EF0100002418";
    attribute INIT_36 of inst : label is "C4089E114E40C199924913AF0000BF25DE91115D4C200764687C90E412952792";
    attribute INIT_37 of inst : label is "0198D109A5459165605554867424AB18D504E34D209105A0785609DE74119584";
    attribute INIT_38 of inst : label is "6C20146768FD4DBAA102645603F9279213F9C0A19564AF034924AF1368395691";
    attribute INIT_39 of inst : label is "65227947AE048931D345225100A10019017576421096E634CC7990B70569115C";
    attribute INIT_3A of inst : label is "10E58D2625C35A55E745552C65267945BF07E140169805F005F055F055F05580";
    attribute INIT_3B of inst : label is "F44975448170951E15E7CB6CCF2C92DF13D46B09159A54E4D450A31991308CDC";
    attribute INIT_3C of inst : label is "9A55E70554E74778B3C95DB2141D50A747596404D65079559C05F6CBA03BCB2C";
    attribute INIT_3D of inst : label is "952B31E4AA00931D3451847F147B11E49D649E64BE0C82CA9331B0C9D8551178";
    attribute INIT_3E of inst : label is "E4248EF7F97A68B06704D3C44323DD02F5C0F510F540F5F0F570A590A5D0A5E0";
    attribute INIT_3F of inst : label is "8193A6DECB684A565AAC2797CF126AA82C661B684A5A623F03C40BC2FD8030E2";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "281E03C01E002D5E3D542D5E07BC003C00782D5E281F3F5502F005F51C2D0B58";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3C0F05783D0C255E";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF0000000000000000333333333333333333333333FFFFFFFF";
    attribute INIT_03 of inst : label is "3333333333333333333333333333333333333333FFFFFFFF2828282807D02D78";
    attribute INIT_04 of inst : label is "3333333333332333333333332333333333333333233333333333333333332233";
    attribute INIT_05 of inst : label is "3333333333333333333333333333333333333333333333333333333333333333";
    attribute INIT_06 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333332D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "3EBCDAA76D229A184C450458489644584845045801F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "76BFFFF7A828FFFF00000000FFE7FEBFFFFFFFFFF82FFFFF0000D007300CDAA7";
    attribute INIT_0D of inst : label is "4281FFFFA96AFC3FA7DAFC3F5FF5F3CF9FF6FD7FE7DBFFFFF96FFFFFFE9FDBFF";
    attribute INIT_0E of inst : label is "7EBD6AA9DEB7F55FE41BFFFFFC3FF28FF3CFF69F3FFCDAA7F82F1FF4AAAAFFFF";
    attribute INIT_0F of inst : label is "E00BFD7FF82FFFFF3FFC6AA9CFF3DAA7F3CFF69FFAAD6BFF6BEBFFE9AFFAF69F";
    attribute INIT_10 of inst : label is "FC3FF41FF00FFFFFDEB7D7D7F7DF2FF807D0C0031FF442817FFD4BE18002F41F";
    attribute INIT_11 of inst : label is "FFFFFFFFAAAAFFFFFC3FFC3FFFFFFFFFFFFFFFFFF6FFFFF656BFFFC1FE9543FF";
    attribute INIT_12 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_14 of inst : label is "AAAA000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "19920510E1E3A91E37A0F415A44FC8A4A93AEA1024501FF901509010FFFF2FF8";
    attribute INIT_16 of inst : label is "F8168291A744DF686386309920100E1E3A91E37A0F015A0E9EAA0A4B3A86386F";
    attribute INIT_17 of inst : label is "AFE638E916FA1A45ABAA4791BA8029EBB278CD0E344A0A6A92AA0AA478CA0790";
    attribute INIT_18 of inst : label is "0F015A838E2A4839ECFBE861F0FE386DB0BEFB3EFA187C3F8E186C2F8E2A4A93";
    attribute INIT_19 of inst : label is "AAA4DE2B0FEEEE1E00CFF03A693A936B1E3790F815A82900E3A25131A479E37A";
    attribute INIT_1A of inst : label is "4A810EB43AD3E6B4FB4FA9ABBBA4DE2A0F0B60BC0EBA1D3E1C3E1C3E1D3E8B9A";
    attribute INIT_1B of inst : label is "E8C0382AE63AE1EF1EF1C71DC71C7BA33032AD8EB9AD3ED4FBBDB00FB53E6D01";
    attribute INIT_1C of inst : label is "935E280F1EF1EF1C71EE8C3EC3EEA2D3ED4FBA00FBA8B4FB4FB071C7B031C71E";
    attribute INIT_1D of inst : label is "AA788AC8EEEEE1E00CF9AFBBAF7BBAFA42FA42F39B41AEC07E1C71DA22E6663D";
    attribute INIT_1E of inst : label is "A91CD2312C43A0AA2928BB58744DD848D6BABA9A9AAABA8AAA9A8A8AAA9ABA8A";
    attribute INIT_1F of inst : label is "786878E5E76A90A0979D59EF224D8A01E67368EA93E83066100103C598401446";
    attribute INIT_20 of inst : label is "3403E00307830082C01CC00BC2D0FA0017350B831F961C9C303830301A340F49";
    attribute INIT_21 of inst : label is "B5001555017A000200545557AD4080000DF80C01017A02AA00E0F81C81F00000";
    attribute INIT_22 of inst : label is "00600C00005A000000C06030A400000002C30E83001F0000C780C2B041000000";
    attribute INIT_23 of inst : label is "00B3038300050000DE00C2C00400000003D00155001E000005C055F0B4000000";
    attribute INIT_24 of inst : label is "00B40055000500001E8057C050000000003500E0000000007800610000000000";
    attribute INIT_25 of inst : label is "002500C0000000005800610000000000003200E300000000F800CB0000000000";
    attribute INIT_26 of inst : label is "0020003300000000A000CC000000000000290015000000006800570000000000";
    attribute INIT_27 of inst : label is "002A000500000000A0005C0000000000002A0018000000008000610000000000";
    attribute INIT_28 of inst : label is "3FFF3FFF015F0000FFFFFFFFFD5000003FFFFFFF07FF00AFFFFCFFFFFFD0FA00";
    attribute INIT_29 of inst : label is "FFFFFFFF057F0000FFFFFFFFFD500000FFFFFFFF057F0000FFFFFFFFFD500000";
    attribute INIT_2A of inst : label is "0B4F039000F8000BF1E006C02F00E000FFFFFFFF057F0000FFFFFFFFFD500000";
    attribute INIT_2B of inst : label is "002F039007F80002F80006C02FD080002FD6F8000015000001E00FFD0D000000";
    attribute INIT_2C of inst : label is "77BFFDEEDFF5FFF024501FF9015090109FD6D8000795000008000FD400000000";
    attribute INIT_2D of inst : label is "341CEFFBCFF3CFF3E7DBDBE7796DB69EF96FDBE7E7DBEFFBDFF7FFFFFEDFFB7F";
    attribute INIT_2E of inst : label is "3FFC3FFCE96BD697D7D7EBEBDBE7E7DBF3CFF3CF7EBDBD7EDFF7382CFFFFFFFF";
    attribute INIT_2F of inst : label is "C7D3CBE3DFF7EFFB3FFC3FFCFC3FFC3FF3CFF3CFFFFC3FFF3FFFFFFCFBEFF7DF";
    attribute INIT_30 of inst : label is "CBE3C7D3D7D7EBEBF82FF41FB7DE7BED20089006382C341C3EBC3D7CC143C283";
    attribute INIT_31 of inst : label is "FFFFFFFFFFFFFFFFCFF3CFF3FFFFFFFFFFFFFFFFF7BFFDEF333FFCCCFCCC333F";
    attribute INIT_32 of inst : label is "AAAAFFFFBBBBAAAABBBBFFFFAAAAEEEEFFFFFFFFAAAABBBBFFFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "00000000AAAAAAAABBBBBBBBEEEEAAAAFFFFBBBBEEEEFFFFEEEEEEEEFFFFAAAA";
    attribute INIT_34 of inst : label is "AAAA555500000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "3C121041A0F2CFC330AC9490C6C2B834CFE38D8D55956A6955559555BFFE7FFD";
    attribute INIT_36 of inst : label is "9882F44CD0C88B3830CB338101840A4F388CC3FA09091F0FEB3B0E4E788F0FB2";
    attribute INIT_37 of inst : label is "E8FB7BB0232E0C4CEFBF3118ACCC3AB3C7BC8B0747974B2FF23B783C2FD3300C";
    attribute INIT_38 of inst : label is "09083C0FCB3B0B30ABA68CF0A2B30FB0A2B3DAAB8F8C0BA2CB0C0BA2CB3B3C0E";
    attribute INIT_39 of inst : label is "B9B8CA3F2E3F8BDE734383F31AA3863A4C2FE22073704CC0E1FB0135C3F0C3FA";
    attribute INIT_3A of inst : label is "694C2C2C2CCBF0BCCFCFAAE2B9F8CA3F1F1E33E03E3F0F730F730F730F73AA0A";
    attribute INIT_3B of inst : label is "F8D04BF687BEB3F63C6DC71C871C78EF50B3EB83BBB03CCCFAFCC383C3B30CC0";
    attribute INIT_3C of inst : label is "D24F0BC33C6DCFD873E78F37B32FB48FCFC38CD8FAEDF3F32D3C71C7C0A1C71E";
    attribute INIT_3D of inst : label is "8FECFF08AAFFB1E53F30FFEADFEAFFAE372E352ECC48E8CC4B9C73C620AA03BD";
    attribute INIT_3E of inst : label is "CEC080691C83E3B74FF0DFDC06C0CE40A73FAFDFAF6FAF9FAF8FAF4FAF9FAFCF";
    attribute INIT_3F of inst : label is "0FB02CB083EBF034F2092E3213CDC80C85EF3BE3E23804A7411061588C045046";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407F8005000F001503C0F";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF05540AAF05501AF5";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFF0000000000000000333333333333333333333333FFFFFFFF";
    attribute INIT_03 of inst : label is "3333333333333333333333333333333333333333FFFFFFFF1414141401400550";
    attribute INIT_04 of inst : label is "3333333333333333333333333333333333333333333333333333333333333333";
    attribute INIT_05 of inst : label is "3333333333333333333333333333333333333333333333333333333333333333";
    attribute INIT_06 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_07 of inst : label is "3333333333333333333333333333333333333333333333331EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "E55B3D7CBC11042C0051472C0071C72C0051472C2ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "EFFFFD6EFFFF7D7F00000000E55BFC3FFFFFFFFFFFFFFD7FE00B0000E55B300C";
    attribute INIT_0D of inst : label is "2FF8F41FFC3F5695FC3F5BE5F3CFAFFAF96FDBE7FEBFF69FFFFFFD7FFFDBF97F";
    attribute INIT_0E of inst : label is "9556BD7EFAAFED7BFFFFD827F14FFC3FF96FF3CFE55B3FFCFFFF8142FFFF5555";
    attribute INIT_0F of inst : label is "FEBFD007FFFFF41F95563FFCE55BCFF3F96FF3CFFFD6B55F97FFD7D6F96F5FF5";
    attribute INIT_10 of inst : label is "F82FFC3FFFFFF00FEBEBED7B1FF4FBEF80020BE081422FF887D2BFFEF82F4001";
    attribute INIT_11 of inst : label is "FFFFFFFFFFFF5555FC3FFC3FFFFFFFFFFFFFFFFF6FFFFF6F83FFFD6AFFC2A97F";
    attribute INIT_12 of inst : label is "0000FFFF00FF000000FFFFFF0000FF00FFFFFFFF000000FFFFFFFFFFFFFFFFFF";
    attribute INIT_13 of inst : label is "000000000000000000FF00FFFF000000FFFF00FFFF00FFFFFF00FF00FFFF0000";
    attribute INIT_14 of inst : label is "0000555500000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0ED010411818F60703C00C50740001D8F60F2D0545555001555515551FF4FFFF";
    attribute INIT_16 of inst : label is "0040F76078400034104100ED010411818B60703C00050747621F1D82C341041C";
    attribute INIT_17 of inst : label is "F03B4076030C1D80EF1D80DC1D800259CF1C030DC73DCB0760F3E1D81C3D03C0";
    attribute INIT_18 of inst : label is "00060743601D80360B0C34100031041C0031C2C30D04000C4104000C401D8F62";
    attribute INIT_19 of inst : label is "00F44B330733331CD2C7303D80C30C30C703C000707C7600D81D831FD83C703C";
    attribute INIT_1A of inst : label is "F10C0D003401CB507507100210F44B3107DC10CC0F531E1F1E1F1E1F1E1F0000";
    attribute INIT_1B of inst : label is "D0F87334073431D41D41C71C071C7343C873400D02D41D4873F0C007C01FBC00";
    attribute INIT_1C of inst : label is "D1CB32071D41D41C71CD0F1F21CF2D41D4873CB873CB5075073C71C7C001C71C";
    attribute INIT_1D of inst : label is "3F2CCCC4333331CD2C7CF4CCD44CCD440D440D4CDC00F300C31C71CC88888B1F";
    attribute INIT_1E of inst : label is "760012012449611F7634DD5C1C005C000F3F3F3F3F2F0F3F2F0F3F2F0F3F1F0F";
    attribute INIT_1F of inst : label is "8C360618180763D060632CB033CF63003D8718476218072B401C701CAD0071C0";
    attribute INIT_20 of inst : label is "D0033803005F0B43C007C02C4100C1E01010373C0111377D1010353505411A96";
    attribute INIT_21 of inst : label is "EAAA6A00000102B5AAA800AD40005E80341F070000000F8180301F8055405E80";
    attribute INIT_22 of inst : label is "0C060300000000250030060000005A000D4301E300000082C170C3400000F800";
    attribute INIT_23 of inst : label is "0343007B00000020C1C0CD000000A0000FAA03A00000002DAA000BC000007800";
    attribute INIT_24 of inst : label is "03AA01780000000AAA002D000000A0000086001E000000000700AE0000000000";
    attribute INIT_25 of inst : label is "0086001A000000000300A4000000000000D3001F00000000C7004C0000000000";
    attribute INIT_26 of inst : label is "0033000500000000CC0004000000000000EA001600000000A800940000000000";
    attribute INIT_27 of inst : label is "003A000500000000A00054000000000000860001000000001800540000000000";
    attribute INIT_28 of inst : label is "3FFF3FFF000002AFFFFFFFFF0000FEA0FFFF3FFF005F0BFFFFFFFFFCF500FFE0";
    attribute INIT_29 of inst : label is "FFFFFFFF00000ABFFFFFFFFF0000FEA0FFFFFFFF00000ABFFFFFFFFF0000FEA0";
    attribute INIT_2A of inst : label is "000001E0001E00BF00000940F400FE00FFFFFFFF00000ABFFFFFFFFF0000FEA0";
    attribute INIT_2B of inst : label is "000009E0006B000B00000B60E900E000F4001FE90000002A0FFE02D000000E00";
    attribute INIT_2C of inst : label is "EFFBDFF7AAAA5FF54555500155551555E4006FE900000B6A0FE8040000000000";
    attribute INIT_2D of inst : label is "6AA9D7D79AA665599EB66D79F7DFFBEF9FF6FD7FFEBFF7DFFBEFDFF7EFDBDBF7";
    attribute INIT_2E of inst : label is "C553CAA3EFFBDFF7EEBBDD77C7D3CBE3DBE7E7DB97D66BE9EBEB9556AAAA5555";
    attribute INIT_2F of inst : label is "EAABD557EBEBD7D795566AA9D697E96BDBE7E7DBE9CBD397F22FF44F9EB66D79";
    attribute INIT_30 of inst : label is "CFF3CFF3EBEBD7D7EFFBDFF77D7DBEBE9416682995566AA9F55FFAAF8AA24551";
    attribute INIT_31 of inst : label is "FFFFFFFFAAAA5555CFF3CFF3FFFFFFFFFFFFFFFF7FFBDFFEE77BDEE7EDDBDBB7";
    attribute INIT_32 of inst : label is "5555FFFF777755557777FFFF5555DDDDFFFFFFFF55557777FFFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "000000005555555577777777DDDD5555FFFF7777DDDDFFFFDDDDDDDDFFFF5555";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "285C04145A05819E244C4D5115816300829E489014101455101400507D7DBEBE";
    attribute INIT_36 of inst : label is "415080B91D8454644104227100102510887952B40405414A06CA380381481341";
    attribute INIT_37 of inst : label is "97A61063165839418A8CE6152840120D9A58470C9668980A20E2A3805A60241C";
    attribute INIT_38 of inst : label is "0407404B0680C0335E195081517013410170E15E48504751041047010600C83B";
    attribute INIT_39 of inst : label is "21204C6B152E4798B10B42F0E0161865855B905006E4008CCA04C25F9E3152B4";
    attribute INIT_3A of inst : label is "C2810D1010D1CD1851C7000721644C68260D63100C1A0F5E0F5A0F5A0F5E0014";
    attribute INIT_3B of inst : label is "F22000E8443871851C51C71D471C40CF88720704214D1F5061FD81438756CC85";
    attribute INIT_3C of inst : label is "B356018B1C51C71473C40F1A73861891F5072AE062CE1471463C71C78051C71C";
    attribute INIT_3D of inst : label is "1AB8B80055AA72841EB1A6959615985058105A1198459488C75872D4BB00CF1B";
    attribute INIT_3E of inst : label is "019C40591681028200AC9A545D4158404E7A0AFA0AEA0A6A0A9A0AAA0A3A0A4A";
    attribute INIT_3F of inst : label is "D86253495C0620C805F779E5338B00897C93580212CC136A0241138598C035C0";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
