library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity splat_prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of splat_prog is
	type rom is array(0 to  49151) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"7E",X"D7",X"AE",X"53",X"50",X"4C",X"41",X"54",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",
		X"49",X"47",X"48",X"54",X"20",X"28",X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",
		X"4C",X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",
		X"43",X"53",X"20",X"49",X"4E",X"43",X"2E",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",
		X"53",X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"8E",X"98",X"24",X"9F",X"1C",X"96",
		X"4B",X"27",X"FC",X"0F",X"4B",X"0C",X"8A",X"D6",X"39",X"2B",X"03",X"7E",X"D1",X"36",X"34",X"01",
		X"1A",X"F0",X"C5",X"40",X"26",X"21",X"96",X"64",X"27",X"1D",X"0A",X"64",X"26",X"19",X"9E",X"66",
		X"27",X"15",X"EC",X"81",X"2B",X"03",X"8E",X"00",X"00",X"9F",X"66",X"D7",X"64",X"C6",X"FF",X"F7",
		X"C8",X"0E",X"84",X"3F",X"B7",X"C8",X"0E",X"35",X"01",X"10",X"8E",X"99",X"6E",X"10",X"9F",X"71",
		X"4F",X"AE",X"A6",X"2A",X"0B",X"BD",X"D7",X"76",X"6F",X"A6",X"8B",X"02",X"81",X"14",X"25",X"F1",
		X"CE",X"00",X"00",X"10",X"8E",X"99",X"BC",X"C6",X"03",X"AE",X"A4",X"27",X"05",X"EF",X"A4",X"BD",
		X"D7",X"84",X"AE",X"22",X"27",X"05",X"EF",X"22",X"BD",X"D7",X"84",X"31",X"A8",X"48",X"5A",X"26",
		X"E8",X"10",X"8E",X"99",X"C0",X"C6",X"03",X"D7",X"3C",X"EC",X"A4",X"27",X"05",X"EF",X"A4",X"BD",
		X"D1",X"5B",X"EC",X"22",X"27",X"05",X"EF",X"22",X"BD",X"D1",X"5B",X"31",X"A8",X"48",X"0A",X"3C",
		X"26",X"E7",X"CE",X"99",X"91",X"C6",X"03",X"D7",X"3C",X"10",X"AE",X"C8",X"33",X"2A",X"05",X"6F",
		X"C8",X"33",X"8D",X"5B",X"10",X"AE",X"C8",X"35",X"2A",X"05",X"6F",X"C8",X"35",X"8D",X"50",X"33",
		X"C8",X"48",X"0A",X"3C",X"26",X"E3",X"BD",X"D3",X"28",X"10",X"8E",X"99",X"91",X"BD",X"D1",X"A3",
		X"10",X"8E",X"99",X"D9",X"BD",X"D1",X"A3",X"10",X"8E",X"9A",X"21",X"BD",X"D1",X"A3",X"BD",X"D4",
		X"38",X"CE",X"99",X"91",X"BD",X"DF",X"0F",X"CE",X"99",X"D9",X"BD",X"DF",X"0F",X"CE",X"9A",X"21",
		X"BD",X"DF",X"0F",X"BD",X"5D",X"BF",X"CE",X"98",X"24",X"20",X"09",X"6A",X"44",X"26",X"05",X"DF",
		X"1C",X"6E",X"D8",X"02",X"EE",X"C4",X"26",X"F3",X"10",X"CE",X"BF",X"00",X"7E",X"D0",X"4A",X"BD",
		X"D6",X"8B",X"5D",X"B3",X"54",X"10",X"AF",X"07",X"EF",X"09",X"39",X"34",X"20",X"1F",X"02",X"8A",
		X"80",X"1F",X"03",X"AE",X"4A",X"AE",X"15",X"A6",X"15",X"8B",X"01",X"A7",X"55",X"A6",X"17",X"A7",
		X"57",X"BD",X"D6",X"8B",X"5D",X"B0",X"22",X"6F",X"09",X"EF",X"07",X"AF",X"4A",X"E6",X"59",X"C4",
		X"0E",X"8E",X"E4",X"F8",X"AE",X"85",X"E6",X"45",X"58",X"58",X"30",X"85",X"EC",X"84",X"10",X"8C",
		X"00",X"00",X"2A",X"04",X"43",X"50",X"82",X"FF",X"ED",X"5C",X"EC",X"02",X"ED",X"5E",X"CE",X"00",
		X"00",X"35",X"A0",X"A6",X"A4",X"10",X"26",X"00",X"82",X"EE",X"3B",X"2B",X"02",X"EE",X"37",X"CC",
		X"25",X"00",X"A3",X"51",X"25",X"35",X"10",X"83",X"06",X"00",X"22",X"04",X"BD",X"D2",X"B1",X"39",
		X"10",X"83",X"26",X"80",X"22",X"F9",X"EE",X"35",X"34",X"20",X"BD",X"D2",X"B1",X"26",X"1A",X"10",
		X"AE",X"E4",X"EE",X"3B",X"2B",X"02",X"EE",X"37",X"BD",X"D2",X"B1",X"26",X"0C",X"10",X"AE",X"E4",
		X"EE",X"3D",X"2B",X"02",X"EE",X"39",X"BD",X"D2",X"B1",X"35",X"A0",X"CC",X"77",X"00",X"A3",X"51",
		X"25",X"09",X"10",X"83",X"06",X"00",X"22",X"04",X"BD",X"D2",X"D2",X"39",X"10",X"83",X"1B",X"00",
		X"22",X"F9",X"EE",X"33",X"2B",X"02",X"EE",X"35",X"34",X"20",X"BD",X"D2",X"D2",X"26",X"1A",X"10",
		X"AE",X"E4",X"EE",X"3B",X"2B",X"02",X"EE",X"37",X"BD",X"D2",X"D2",X"26",X"0C",X"10",X"AE",X"E4",
		X"EE",X"3D",X"2B",X"02",X"EE",X"39",X"BD",X"D2",X"D2",X"35",X"A0",X"EE",X"3D",X"2B",X"02",X"EE",
		X"39",X"EC",X"51",X"83",X"6A",X"00",X"25",X"39",X"10",X"83",X"06",X"00",X"22",X"04",X"BD",X"D2",
		X"D2",X"39",X"10",X"83",X"1B",X"00",X"22",X"F9",X"EE",X"33",X"2B",X"02",X"EE",X"35",X"34",X"20",
		X"BD",X"D2",X"D2",X"26",X"1A",X"10",X"AE",X"E4",X"EE",X"3D",X"2B",X"02",X"EE",X"39",X"BD",X"D2",
		X"D2",X"26",X"0C",X"10",X"AE",X"E4",X"EE",X"3B",X"2B",X"02",X"EE",X"37",X"BD",X"D2",X"D2",X"35",
		X"A0",X"EC",X"51",X"83",X"18",X"00",X"25",X"09",X"10",X"83",X"06",X"00",X"22",X"04",X"BD",X"D2",
		X"B1",X"39",X"10",X"83",X"1B",X"00",X"22",X"F9",X"EE",X"33",X"2B",X"02",X"EE",X"35",X"34",X"20",
		X"BD",X"D2",X"B1",X"26",X"1A",X"10",X"AE",X"E4",X"EE",X"3D",X"2B",X"02",X"EE",X"39",X"BD",X"D2",
		X"B1",X"26",X"0C",X"10",X"AE",X"E4",X"EE",X"3B",X"2B",X"02",X"EE",X"37",X"BD",X"D2",X"B1",X"35",
		X"A0",X"A6",X"53",X"9E",X"6B",X"9C",X"69",X"27",X"17",X"8C",X"99",X"1E",X"26",X"03",X"8E",X"99",
		X"46",X"10",X"AE",X"83",X"27",X"EF",X"A1",X"34",X"22",X"EB",X"E6",X"54",X"E1",X"33",X"24",X"23",
		X"5F",X"39",X"A6",X"53",X"9E",X"6F",X"9C",X"6D",X"27",X"17",X"8C",X"99",X"46",X"26",X"03",X"8E",
		X"99",X"6E",X"10",X"AE",X"83",X"27",X"EF",X"A1",X"34",X"22",X"EB",X"E6",X"54",X"E1",X"33",X"22",
		X"02",X"5F",X"39",X"A6",X"33",X"A1",X"53",X"23",X"06",X"30",X"C4",X"33",X"A4",X"20",X"02",X"30",
		X"A4",X"EC",X"11",X"10",X"A3",X"51",X"23",X"10",X"10",X"AE",X"5A",X"EC",X"51",X"AB",X"3E",X"10",
		X"A3",X"11",X"10",X"22",X"00",X"A7",X"5F",X"39",X"10",X"AE",X"1A",X"EC",X"11",X"AB",X"3E",X"10",
		X"A3",X"51",X"10",X"22",X"00",X"BD",X"20",X"EE",X"8E",X"98",X"2A",X"9F",X"60",X"AE",X"84",X"10",
		X"27",X"00",X"7B",X"EE",X"84",X"27",X"26",X"A6",X"13",X"A1",X"53",X"22",X"06",X"9F",X"60",X"AE",
		X"84",X"20",X"F0",X"DF",X"62",X"EE",X"C4",X"27",X"04",X"A1",X"53",X"22",X"F6",X"10",X"AE",X"84",
		X"10",X"AF",X"9F",X"98",X"60",X"EF",X"84",X"AF",X"9F",X"98",X"62",X"20",X"CB",X"8E",X"98",X"2A",
		X"20",X"46",X"A6",X"14",X"A1",X"53",X"25",X"40",X"E6",X"03",X"27",X"04",X"E5",X"43",X"26",X"34",
		X"E6",X"11",X"27",X"34",X"A6",X"51",X"27",X"2C",X"E1",X"51",X"25",X"15",X"10",X"AE",X"5A",X"AB",
		X"3E",X"E6",X"52",X"2A",X"06",X"A1",X"11",X"25",X"1B",X"20",X"24",X"A1",X"11",X"23",X"15",X"20",
		X"1E",X"10",X"AE",X"1A",X"EB",X"3E",X"A6",X"12",X"2A",X"06",X"E1",X"51",X"25",X"06",X"20",X"16",
		X"E1",X"51",X"22",X"12",X"EE",X"C4",X"26",X"BA",X"AE",X"84",X"EE",X"84",X"26",X"B4",X"39",X"CC",
		X"D3",X"A4",X"34",X"06",X"20",X"07",X"CC",X"D3",X"A4",X"34",X"06",X"20",X"26",X"BD",X"D4",X"16",
		X"31",X"21",X"A6",X"A4",X"2B",X"4C",X"44",X"56",X"C4",X"80",X"E3",X"51",X"DD",X"43",X"A6",X"84",
		X"2B",X"40",X"44",X"56",X"C4",X"80",X"D3",X"3F",X"10",X"93",X"43",X"23",X"2C",X"30",X"02",X"31",
		X"22",X"20",X"DF",X"BD",X"D4",X"16",X"30",X"01",X"A6",X"A4",X"2B",X"26",X"44",X"56",X"C4",X"80",
		X"E3",X"51",X"DD",X"43",X"A6",X"84",X"2B",X"1A",X"44",X"56",X"C4",X"80",X"D3",X"3F",X"10",X"93",
		X"43",X"24",X"06",X"30",X"02",X"31",X"22",X"20",X"DF",X"9E",X"41",X"AF",X"46",X"EF",X"06",X"C6",
		X"01",X"39",X"9E",X"41",X"5F",X"39",X"A6",X"53",X"A0",X"13",X"97",X"3C",X"EC",X"11",X"DD",X"3F",
		X"9F",X"41",X"10",X"AE",X"1A",X"EC",X"3E",X"3D",X"30",X"AB",X"96",X"3C",X"48",X"30",X"86",X"10",
		X"AE",X"5A",X"EC",X"3E",X"3D",X"31",X"AB",X"39",X"10",X"9E",X"69",X"10",X"9C",X"6B",X"27",X"1A",
		X"AE",X"A1",X"27",X"09",X"A6",X"11",X"26",X"12",X"BD",X"D7",X"76",X"0C",X"90",X"10",X"8C",X"99",
		X"46",X"26",X"04",X"10",X"8E",X"99",X"1E",X"10",X"9F",X"69",X"10",X"9E",X"6D",X"10",X"9C",X"6F",
		X"27",X"1A",X"AE",X"A1",X"27",X"09",X"A6",X"11",X"26",X"12",X"BD",X"D7",X"76",X"0C",X"91",X"10",
		X"8C",X"99",X"6E",X"26",X"04",X"10",X"8E",X"99",X"46",X"10",X"9F",X"6D",X"10",X"9E",X"69",X"10",
		X"9C",X"6B",X"27",X"3F",X"AE",X"A1",X"27",X"2F",X"5F",X"A6",X"11",X"10",X"83",X"1E",X"00",X"23",
		X"19",X"9F",X"3F",X"AE",X"1A",X"A6",X"1E",X"9E",X"3F",X"AB",X"11",X"10",X"83",X"2A",X"00",X"22",
		X"10",X"EC",X"1E",X"C3",X"00",X"06",X"ED",X"1E",X"20",X"07",X"86",X"01",X"ED",X"1E",X"4F",X"ED",
		X"1C",X"A6",X"06",X"27",X"02",X"8D",X"4B",X"10",X"8C",X"99",X"46",X"26",X"C2",X"10",X"8E",X"99",
		X"1E",X"20",X"BC",X"10",X"9E",X"6D",X"10",X"9C",X"6F",X"10",X"27",X"01",X"0A",X"AE",X"A1",X"27",
		X"25",X"EC",X"11",X"5F",X"10",X"83",X"70",X"00",X"24",X"0F",X"10",X"83",X"6B",X"00",X"25",X"10",
		X"EC",X"1E",X"C3",X"00",X"06",X"ED",X"1E",X"20",X"07",X"86",X"01",X"ED",X"1E",X"4F",X"ED",X"1C",
		X"A6",X"06",X"27",X"02",X"8D",X"0C",X"10",X"8C",X"99",X"6E",X"26",X"CA",X"10",X"8E",X"99",X"46",
		X"20",X"C4",X"10",X"9F",X"43",X"EE",X"06",X"A6",X"59",X"85",X"C0",X"26",X"18",X"10",X"9E",X"43",
		X"CC",X"00",X"00",X"ED",X"3E",X"1A",X"50",X"6F",X"15",X"DE",X"71",X"AF",X"C1",X"DF",X"71",X"BD",
		X"DC",X"73",X"1C",X"AF",X"39",X"10",X"AE",X"4A",X"85",X"40",X"27",X"15",X"4F",X"E6",X"11",X"E1",
		X"51",X"22",X"04",X"E6",X"3B",X"27",X"0A",X"4C",X"E6",X"3D",X"2A",X"05",X"4A",X"E6",X"3B",X"26",
		X"CC",X"E6",X"33",X"27",X"0F",X"BD",X"D7",X"20",X"BD",X"D5",X"5A",X"10",X"9E",X"43",X"CC",X"00",
		X"00",X"ED",X"3E",X"39",X"6F",X"06",X"10",X"9E",X"43",X"39",X"34",X"41",X"5F",X"E7",X"06",X"6C",
		X"02",X"BD",X"DC",X"73",X"10",X"AE",X"4A",X"10",X"AF",X"0A",X"85",X"01",X"27",X"33",X"A6",X"19",
		X"85",X"01",X"26",X"06",X"8A",X"01",X"A7",X"19",X"8D",X"47",X"4F",X"A7",X"46",X"ED",X"1C",X"ED",
		X"1E",X"1A",X"50",X"AF",X"3D",X"AE",X"39",X"A6",X"03",X"10",X"AE",X"3D",X"A7",X"23",X"A6",X"04",
		X"A7",X"25",X"BD",X"D8",X"D8",X"6F",X"22",X"EC",X"35",X"ED",X"31",X"A6",X"37",X"A7",X"33",X"35",
		X"C1",X"A6",X"19",X"85",X"01",X"27",X"06",X"84",X"0E",X"A7",X"19",X"8D",X"14",X"4F",X"A7",X"46",
		X"ED",X"1C",X"ED",X"1E",X"1A",X"50",X"AF",X"3B",X"AE",X"37",X"A6",X"03",X"10",X"AE",X"3B",X"20",
		X"CB",X"34",X"24",X"10",X"8E",X"00",X"00",X"48",X"10",X"AE",X"A6",X"10",X"AF",X"08",X"EC",X"A4",
		X"C3",X"00",X"02",X"ED",X"1A",X"35",X"A4",X"96",X"68",X"27",X"3D",X"0A",X"68",X"26",X"39",X"B6",
		X"99",X"04",X"97",X"68",X"8D",X"33",X"86",X"3D",X"A0",X"5E",X"10",X"8E",X"FF",X"D0",X"8D",X"71",
		X"DE",X"6B",X"AF",X"C1",X"11",X"83",X"99",X"46",X"26",X"03",X"CE",X"99",X"1E",X"DF",X"6B",X"8D",
		X"18",X"86",X"58",X"10",X"8E",X"00",X"30",X"8D",X"58",X"DE",X"6F",X"AF",X"C1",X"11",X"83",X"99",
		X"6E",X"26",X"03",X"CE",X"99",X"46",X"DF",X"6F",X"39",X"9E",X"30",X"26",X"01",X"3F",X"EC",X"84",
		X"DD",X"30",X"DC",X"2C",X"ED",X"84",X"CE",X"D4",X"38",X"EF",X"0A",X"6F",X"06",X"6F",X"0C",X"6F",
		X"03",X"BD",X"5D",X"BF",X"4A",X"90",X"BA",X"86",X"05",X"25",X"0A",X"96",X"73",X"2A",X"06",X"BD",
		X"5D",X"BF",X"C6",X"05",X"3D",X"48",X"A7",X"19",X"48",X"CE",X"00",X"00",X"EE",X"C6",X"EF",X"08",
		X"EE",X"C4",X"C6",X"2B",X"E7",X"14",X"E0",X"41",X"E7",X"17",X"E7",X"13",X"33",X"42",X"EF",X"1A",
		X"39",X"5F",X"ED",X"11",X"ED",X"15",X"4F",X"5F",X"ED",X"1E",X"A7",X"18",X"A7",X"04",X"A7",X"05",
		X"10",X"AF",X"1C",X"9F",X"2C",X"39",X"34",X"62",X"DE",X"28",X"26",X"01",X"3F",X"10",X"AE",X"C4",
		X"10",X"9F",X"28",X"86",X"01",X"A7",X"46",X"A6",X"E4",X"20",X"19",X"35",X"10",X"30",X"03",X"34",
		X"10",X"A6",X"1F",X"AE",X"1D",X"34",X"62",X"DE",X"26",X"26",X"01",X"3F",X"10",X"AE",X"C4",X"10",
		X"9F",X"26",X"6F",X"46",X"AF",X"42",X"A7",X"45",X"86",X"01",X"A7",X"44",X"AE",X"9F",X"98",X"1C",
		X"EF",X"9F",X"98",X"1C",X"AF",X"C4",X"30",X"C4",X"35",X"E2",X"AE",X"E1",X"DE",X"1C",X"A7",X"44",
		X"AF",X"42",X"7E",X"D1",X"44",X"9E",X"1C",X"8D",X"07",X"33",X"84",X"7E",X"D1",X"44",X"AE",X"0A",
		X"34",X"46",X"CE",X"98",X"24",X"AC",X"C4",X"26",X"18",X"EC",X"84",X"ED",X"C4",X"A6",X"06",X"27",
		X"06",X"DC",X"28",X"9F",X"28",X"20",X"04",X"DC",X"26",X"9F",X"26",X"ED",X"84",X"30",X"C4",X"35",
		X"C6",X"EE",X"C4",X"26",X"E0",X"3F",X"34",X"10",X"8E",X"98",X"24",X"20",X"0A",X"A1",X"05",X"26",
		X"06",X"9C",X"1C",X"27",X"02",X"8D",X"C9",X"AE",X"84",X"26",X"F2",X"35",X"90",X"34",X"12",X"8E",
		X"98",X"24",X"20",X"06",X"9C",X"1C",X"27",X"02",X"8D",X"B6",X"AE",X"84",X"26",X"F6",X"35",X"92",
		X"34",X"46",X"CE",X"98",X"2C",X"AC",X"C4",X"26",X"0E",X"EC",X"D4",X"ED",X"C4",X"DC",X"2A",X"9F",
		X"2A",X"ED",X"84",X"6F",X"02",X"35",X"C6",X"EE",X"C4",X"26",X"EA",X"3F",X"8D",X"12",X"34",X"46",
		X"EF",X"0A",X"EE",X"64",X"37",X"06",X"ED",X"08",X"37",X"02",X"A7",X"03",X"EF",X"64",X"35",X"C6",
		X"34",X"06",X"9E",X"30",X"26",X"01",X"3F",X"EC",X"84",X"DD",X"30",X"DC",X"2A",X"ED",X"84",X"CC",
		X"00",X"00",X"ED",X"11",X"A7",X"13",X"ED",X"1C",X"ED",X"1E",X"A7",X"19",X"A7",X"06",X"A7",X"02",
		X"ED",X"04",X"A7",X"0C",X"35",X"86",X"34",X"56",X"CE",X"98",X"2C",X"20",X"0C",X"34",X"56",X"CE",
		X"98",X"2E",X"20",X"05",X"34",X"56",X"CE",X"98",X"2A",X"AC",X"C4",X"26",X"0C",X"EC",X"D4",X"ED",
		X"C4",X"DC",X"30",X"9F",X"30",X"ED",X"84",X"35",X"D6",X"EE",X"C4",X"26",X"EC",X"3F",X"00",X"34",
		X"FF",X"35",X"00",X"34",X"00",X"3E",X"C8",X"0C",X"C8",X"0E",X"C8",X"04",X"C8",X"06",X"1A",X"FF",
		X"10",X"CE",X"BF",X"00",X"86",X"98",X"1F",X"8B",X"86",X"01",X"B7",X"C9",X"00",X"8E",X"D7",X"9E",
		X"4F",X"5F",X"ED",X"98",X"08",X"EC",X"81",X"ED",X"98",X"06",X"8C",X"D7",X"A6",X"26",X"F1",X"86",
		X"FF",X"B7",X"C8",X"0E",X"86",X"3F",X"B7",X"C8",X"0E",X"BD",X"DD",X"0F",X"8E",X"98",X"00",X"C6",
		X"39",X"6F",X"80",X"F7",X"CB",X"FF",X"8C",X"BF",X"7F",X"26",X"F6",X"CC",X"A5",X"5A",X"DD",X"20",
		X"CC",X"70",X"FF",X"DD",X"35",X"CC",X"0E",X"10",X"DD",X"49",X"8E",X"CD",X"00",X"BD",X"37",X"C2",
		X"1F",X"98",X"81",X"20",X"22",X"06",X"84",X"0F",X"81",X"09",X"23",X"07",X"5F",X"8E",X"CD",X"00",
		X"BD",X"37",X"CB",X"F7",X"BF",X"32",X"8D",X"14",X"8D",X"53",X"8D",X"40",X"BD",X"D8",X"F1",X"BD",
		X"D6",X"8B",X"5D",X"A7",X"31",X"0F",X"1E",X"1C",X"00",X"7E",X"D0",X"4A",X"34",X"16",X"CC",X"00",
		X"00",X"8E",X"A2",X"8E",X"9F",X"26",X"30",X"0F",X"AF",X"11",X"8C",X"A5",X"6D",X"26",X"F7",X"ED",
		X"84",X"DD",X"24",X"8E",X"A5",X"7C",X"9F",X"28",X"30",X"88",X"44",X"AF",X"88",X"BC",X"8C",X"AA",
		X"88",X"26",X"F5",X"ED",X"84",X"8E",X"98",X"24",X"9F",X"1C",X"35",X"96",X"8E",X"DD",X"2F",X"CE",
		X"98",X"00",X"EC",X"81",X"ED",X"C1",X"11",X"83",X"98",X"10",X"25",X"F6",X"39",X"34",X"17",X"1A",
		X"50",X"8E",X"9A",X"69",X"9F",X"30",X"30",X"88",X"1C",X"AF",X"88",X"E4",X"8C",X"A2",X"81",X"26",
		X"F5",X"CC",X"00",X"00",X"ED",X"84",X"DD",X"2C",X"DD",X"2A",X"DD",X"2E",X"35",X"97",X"1F",X"20",
		X"5F",X"ED",X"11",X"ED",X"15",X"1F",X"20",X"E7",X"13",X"8D",X"2B",X"1F",X"98",X"5F",X"ED",X"17",
		X"E7",X"04",X"E7",X"05",X"86",X"40",X"A7",X"19",X"9F",X"2A",X"39",X"8E",X"98",X"3A",X"C6",X"39",
		X"4F",X"A7",X"80",X"F7",X"CB",X"FF",X"8C",X"9A",X"5A",X"26",X"F6",X"86",X"FF",X"B7",X"C8",X"0E",
		X"86",X"1F",X"B7",X"C8",X"0E",X"39",X"34",X"44",X"E6",X"13",X"EE",X"08",X"EE",X"C4",X"EB",X"41",
		X"E7",X"14",X"33",X"42",X"EF",X"1A",X"35",X"C4",X"34",X"46",X"EE",X"28",X"86",X"05",X"E6",X"25",
		X"3D",X"33",X"C5",X"EC",X"42",X"E3",X"15",X"ED",X"35",X"A6",X"44",X"AB",X"17",X"A7",X"37",X"35",
		X"C6",X"CC",X"99",X"1E",X"DD",X"69",X"DD",X"6B",X"CC",X"99",X"46",X"DD",X"6D",X"DD",X"6F",X"86",
		X"0F",X"97",X"68",X"39",X"34",X"04",X"5F",X"81",X"10",X"25",X"06",X"CB",X"0A",X"80",X"10",X"20",
		X"F6",X"34",X"04",X"AB",X"E0",X"35",X"84",X"34",X"04",X"1F",X"89",X"4F",X"C1",X"0A",X"25",X"07",
		X"8B",X"10",X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",X"AB",X"E0",X"19",X"35",X"84",X"86",X"98",
		X"1F",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"86",X"34",X"B7",X"C8",X"0F",X"B6",X"C8",X"0E",X"B6",
		X"CB",X"00",X"97",X"5E",X"10",X"2B",X"00",X"D3",X"81",X"06",X"22",X"1B",X"CE",X"C0",X"10",X"DC",
		X"0A",X"9E",X"0C",X"10",X"9E",X"0E",X"36",X"36",X"DC",X"04",X"9E",X"06",X"10",X"9E",X"08",X"36",
		X"36",X"DC",X"00",X"9E",X"02",X"36",X"16",X"B6",X"CB",X"00",X"84",X"C0",X"10",X"26",X"00",X"9B",
		X"96",X"39",X"2A",X"14",X"48",X"2B",X"11",X"DC",X"49",X"83",X"00",X"01",X"2E",X"08",X"C6",X"06",
		X"BD",X"37",X"B9",X"CC",X"0E",X"10",X"DD",X"49",X"96",X"12",X"27",X"02",X"0A",X"12",X"DC",X"19",
		X"DD",X"1A",X"DC",X"17",X"DD",X"18",X"DC",X"15",X"DD",X"16",X"DC",X"13",X"DD",X"14",X"B6",X"C8",
		X"0C",X"97",X"13",X"85",X"40",X"27",X"04",X"C6",X"78",X"D7",X"12",X"D6",X"13",X"DA",X"14",X"DA",
		X"15",X"DA",X"16",X"DA",X"17",X"DA",X"18",X"DA",X"19",X"DA",X"1A",X"DA",X"1B",X"D4",X"10",X"D7",
		X"11",X"94",X"14",X"9A",X"11",X"D6",X"10",X"97",X"10",X"53",X"1F",X"98",X"D4",X"10",X"C4",X"0A",
		X"9A",X"10",X"43",X"84",X"34",X"A7",X"E2",X"EA",X"E4",X"54",X"27",X"2D",X"E7",X"E4",X"64",X"E4",
		X"24",X"03",X"BD",X"F0",X"03",X"64",X"E4",X"24",X"07",X"96",X"12",X"26",X"03",X"BD",X"37",X"DA",
		X"64",X"E4",X"24",X"03",X"BD",X"37",X"B3",X"96",X"12",X"26",X"0E",X"64",X"E4",X"24",X"03",X"BD",
		X"37",X"D4",X"64",X"E4",X"24",X"03",X"BD",X"37",X"D7",X"35",X"04",X"BD",X"DA",X"4B",X"0D",X"1E",
		X"27",X"2C",X"0F",X"1E",X"DC",X"36",X"BD",X"DA",X"B1",X"20",X"23",X"BD",X"DA",X"4B",X"0D",X"1E",
		X"26",X"1C",X"0C",X"1E",X"0C",X"4B",X"BD",X"5D",X"AA",X"BD",X"DA",X"91",X"B6",X"CB",X"00",X"80",
		X"17",X"81",X"D0",X"23",X"02",X"86",X"D0",X"97",X"37",X"DC",X"37",X"BD",X"DA",X"B1",X"7D",X"C8",
		X"0F",X"10",X"2B",X"FE",X"E9",X"86",X"35",X"B7",X"C8",X"0F",X"3B",X"C6",X"3C",X"F7",X"C8",X"07",
		X"8E",X"99",X"91",X"CE",X"98",X"56",X"8D",X"0A",X"8E",X"99",X"D9",X"33",X"44",X"86",X"34",X"B7",
		X"C8",X"07",X"B6",X"C8",X"04",X"34",X"02",X"A4",X"C4",X"AA",X"42",X"A7",X"42",X"A6",X"E4",X"AA",
		X"C4",X"A4",X"42",X"A7",X"42",X"35",X"02",X"A7",X"C4",X"B6",X"C8",X"06",X"34",X"02",X"A4",X"41",
		X"AA",X"43",X"A7",X"43",X"A6",X"E4",X"AA",X"41",X"A4",X"43",X"A7",X"43",X"35",X"02",X"A7",X"41",
		X"39",X"8E",X"98",X"2C",X"8D",X"16",X"8E",X"98",X"2A",X"8D",X"11",X"8E",X"98",X"2E",X"20",X"0C",
		X"EC",X"15",X"E3",X"1C",X"ED",X"15",X"EC",X"17",X"E3",X"1E",X"ED",X"17",X"AE",X"84",X"26",X"F0",
		X"39",X"DD",X"34",X"8E",X"98",X"2C",X"0F",X"3A",X"0F",X"4D",X"BD",X"DB",X"F9",X"86",X"08",X"97",
		X"4D",X"96",X"39",X"10",X"2A",X"00",X"BA",X"CE",X"99",X"91",X"AE",X"53",X"2B",X"0C",X"AE",X"55",
		X"96",X"5F",X"80",X"04",X"97",X"5F",X"2A",X"02",X"0C",X"3A",X"A6",X"17",X"91",X"34",X"10",X"22",
		X"00",X"92",X"91",X"35",X"10",X"25",X"00",X"8C",X"E6",X"02",X"10",X"26",X"00",X"86",X"AE",X"55",
		X"BD",X"DC",X"73",X"AE",X"59",X"BD",X"DC",X"73",X"AE",X"57",X"BD",X"DC",X"73",X"AE",X"5D",X"2A",
		X"03",X"BD",X"DC",X"73",X"AE",X"5B",X"2A",X"03",X"BD",X"DC",X"73",X"AE",X"53",X"2A",X"03",X"BD",
		X"DC",X"73",X"DF",X"4E",X"AE",X"55",X"E6",X"11",X"27",X"09",X"E6",X"02",X"26",X"05",X"BD",X"DC",
		X"A0",X"DE",X"4E",X"AE",X"59",X"E6",X"11",X"27",X"09",X"E6",X"02",X"26",X"05",X"BD",X"DC",X"A0",
		X"DE",X"4E",X"AE",X"57",X"E6",X"11",X"27",X"09",X"E6",X"02",X"26",X"05",X"BD",X"DC",X"A0",X"DE",
		X"4E",X"AE",X"5D",X"2A",X"0D",X"E6",X"11",X"27",X"09",X"E6",X"02",X"26",X"05",X"BD",X"DC",X"A0",
		X"DE",X"4E",X"AE",X"5B",X"2A",X"0D",X"E6",X"11",X"27",X"09",X"E6",X"02",X"26",X"05",X"BD",X"DC",
		X"A0",X"DE",X"4E",X"AE",X"53",X"2A",X"0D",X"E6",X"11",X"27",X"09",X"E6",X"02",X"26",X"05",X"BD",
		X"DC",X"A0",X"DE",X"4E",X"0F",X"3A",X"33",X"C8",X"48",X"11",X"83",X"9A",X"21",X"10",X"23",X"FF",
		X"49",X"8E",X"98",X"2A",X"8D",X"53",X"8E",X"98",X"2E",X"0C",X"3A",X"8D",X"4C",X"7E",X"DB",X"FE",
		X"E6",X"0A",X"C1",X"9A",X"22",X"07",X"EE",X"0A",X"AC",X"C8",X"27",X"26",X"3C",X"A6",X"17",X"91",
		X"34",X"22",X"36",X"91",X"35",X"25",X"32",X"A6",X"11",X"27",X"2E",X"E6",X"02",X"26",X"2A",X"EE",
		X"1A",X"E6",X"13",X"FD",X"CA",X"04",X"EC",X"5E",X"FD",X"CA",X"06",X"FF",X"CA",X"02",X"7F",X"CA",
		X"01",X"C6",X"1A",X"6D",X"12",X"2A",X"02",X"CA",X"20",X"F7",X"CA",X"00",X"A6",X"15",X"26",X"06",
		X"A7",X"11",X"A7",X"12",X"20",X"03",X"BD",X"DC",X"A0",X"AE",X"84",X"26",X"B3",X"39",X"A6",X"17",
		X"91",X"34",X"22",X"15",X"91",X"35",X"25",X"11",X"A6",X"11",X"27",X"0D",X"A6",X"15",X"26",X"06",
		X"A7",X"11",X"A7",X"12",X"20",X"03",X"BD",X"DC",X"9A",X"AE",X"84",X"26",X"E1",X"39",X"96",X"39",
		X"2A",X"48",X"96",X"5E",X"2A",X"0B",X"86",X"01",X"8D",X"0C",X"4C",X"8D",X"09",X"86",X"04",X"20",
		X"05",X"4F",X"8D",X"02",X"86",X"03",X"8E",X"98",X"AD",X"E6",X"86",X"2B",X"2D",X"34",X"04",X"8E",
		X"98",X"B2",X"E1",X"86",X"27",X"07",X"7F",X"CA",X"01",X"C6",X"1A",X"8D",X"1E",X"35",X"04",X"E7",
		X"86",X"8E",X"98",X"A8",X"E6",X"86",X"F7",X"CA",X"01",X"27",X"04",X"C6",X"1A",X"20",X"02",X"C6",
		X"0A",X"8E",X"98",X"AD",X"8D",X"05",X"C6",X"FF",X"E7",X"86",X"39",X"34",X"46",X"A6",X"86",X"C6",
		X"14",X"3D",X"C3",X"E9",X"36",X"1F",X"03",X"A6",X"E4",X"48",X"48",X"33",X"C6",X"EC",X"42",X"FD",
		X"CA",X"04",X"EE",X"C4",X"EC",X"C1",X"FD",X"CA",X"06",X"FF",X"CA",X"02",X"A6",X"61",X"B7",X"CA",
		X"00",X"35",X"C6",X"34",X"47",X"1A",X"50",X"EE",X"1A",X"A6",X"11",X"27",X"1B",X"E6",X"13",X"FD",
		X"CA",X"04",X"EC",X"5E",X"FD",X"CA",X"06",X"FF",X"CA",X"02",X"7F",X"CA",X"01",X"C6",X"1A",X"A6",
		X"12",X"2A",X"02",X"CA",X"20",X"F7",X"CA",X"00",X"35",X"C7",X"E6",X"17",X"A6",X"15",X"20",X"0C",
		X"A6",X"15",X"81",X"06",X"25",X"57",X"E6",X"17",X"C1",X"37",X"25",X"51",X"E7",X"13",X"FD",X"CA",
		X"04",X"A7",X"11",X"A6",X"05",X"A1",X"04",X"27",X"0F",X"A7",X"04",X"C6",X"05",X"3D",X"EE",X"08",
		X"EE",X"C5",X"33",X"42",X"EF",X"1A",X"20",X"02",X"EE",X"1A",X"EC",X"5E",X"FD",X"CA",X"06",X"EB",
		X"13",X"E7",X"14",X"C1",X"E7",X"22",X"26",X"AB",X"11",X"81",X"90",X"22",X"20",X"FF",X"CA",X"02",
		X"86",X"02",X"9A",X"4D",X"E6",X"16",X"2A",X"02",X"8A",X"20",X"E7",X"12",X"D6",X"3A",X"27",X"09",
		X"E6",X"0C",X"27",X"05",X"F7",X"CA",X"01",X"8A",X"10",X"B7",X"CA",X"00",X"39",X"96",X"4D",X"26",
		X"09",X"EC",X"17",X"A3",X"1E",X"A7",X"13",X"BD",X"DC",X"73",X"6F",X"11",X"6F",X"12",X"39",X"34",
		X"76",X"CE",X"98",X"00",X"8E",X"00",X"00",X"1F",X"12",X"1F",X"10",X"36",X"36",X"36",X"36",X"36",
		X"36",X"36",X"36",X"36",X"36",X"36",X"10",X"11",X"83",X"00",X"00",X"26",X"EE",X"35",X"F6",X"00",
		X"FF",X"2F",X"5F",X"0F",X"18",X"E0",X"0C",X"D0",X"16",X"4A",X"52",X"04",X"9C",X"02",X"80",X"86",
		X"2C",X"A7",X"49",X"6F",X"48",X"6F",X"47",X"96",X"8B",X"BD",X"D6",X"BA",X"8E",X"94",X"1D",X"A6",
		X"48",X"85",X"02",X"27",X"04",X"30",X"89",X"FF",X"00",X"81",X"01",X"27",X"06",X"81",X"02",X"27",
		X"02",X"30",X"1F",X"10",X"8E",X"DD",X"FC",X"BD",X"DD",X"D5",X"A6",X"47",X"44",X"E6",X"A6",X"25",
		X"04",X"54",X"54",X"54",X"54",X"C4",X"0F",X"27",X"2A",X"A6",X"48",X"97",X"3C",X"1F",X"98",X"84",
		X"03",X"54",X"54",X"04",X"3C",X"25",X"07",X"1E",X"89",X"04",X"3C",X"25",X"06",X"50",X"04",X"3C",
		X"24",X"02",X"50",X"40",X"9F",X"3F",X"9B",X"3F",X"DB",X"40",X"1F",X"01",X"BD",X"DD",X"D5",X"6C",
		X"47",X"20",X"C7",X"A6",X"47",X"81",X"69",X"27",X"04",X"6C",X"47",X"20",X"0C",X"6F",X"47",X"6C",
		X"48",X"A6",X"48",X"81",X"04",X"26",X"02",X"6F",X"48",X"6A",X"49",X"10",X"26",X"FF",X"88",X"4F",
		X"97",X"75",X"97",X"86",X"97",X"85",X"4C",X"97",X"D1",X"97",X"C9",X"86",X"07",X"BD",X"D6",X"BA",
		X"0A",X"8D",X"7E",X"D6",X"C5",X"34",X"21",X"1A",X"50",X"7F",X"C9",X"00",X"1F",X"10",X"44",X"1F",
		X"02",X"1F",X"10",X"E6",X"A4",X"85",X"01",X"26",X"06",X"C4",X"0F",X"DA",X"8F",X"20",X"04",X"C4",
		X"F0",X"DA",X"8E",X"E7",X"A4",X"86",X"01",X"B7",X"C9",X"00",X"35",X"A1",X"11",X"11",X"11",X"11",
		X"10",X"33",X"51",X"10",X"35",X"11",X"51",X"14",X"06",X"15",X"11",X"41",X"14",X"14",X"06",X"55",
		X"14",X"11",X"41",X"40",X"55",X"55",X"41",X"14",X"14",X"0E",X"54",X"51",X"41",X"40",X"94",X"54",
		X"55",X"41",X"40",X"98",X"44",X"14",X"14",X"41",X"04",X"4D",X"84",X"14",X"0C",X"44",X"44",X"44",
		X"10",X"34",X"02",X"86",X"01",X"58",X"26",X"04",X"E6",X"C0",X"58",X"5C",X"49",X"6A",X"E4",X"26",
		X"F4",X"32",X"61",X"39",X"8E",X"00",X"30",X"10",X"8E",X"00",X"20",X"CE",X"23",X"BB",X"34",X"16",
		X"6F",X"E4",X"E6",X"E4",X"4F",X"4C",X"58",X"26",X"04",X"E6",X"C0",X"58",X"5C",X"24",X"F6",X"8D",
		X"D0",X"80",X"02",X"A7",X"61",X"86",X"03",X"8D",X"C8",X"E7",X"E4",X"E6",X"61",X"26",X"35",X"84",
		X"07",X"27",X"2F",X"0D",X"39",X"2B",X"25",X"9E",X"1C",X"10",X"AF",X"08",X"EF",X"07",X"35",X"66",
		X"A7",X"0A",X"10",X"AF",X"0B",X"EF",X"0D",X"86",X"01",X"BD",X"D6",X"BA",X"10",X"AE",X"4D",X"AE",
		X"4B",X"A6",X"4A",X"34",X"36",X"E6",X"49",X"4F",X"1F",X"02",X"EE",X"47",X"AE",X"62",X"31",X"21",
		X"20",X"B0",X"35",X"96",X"84",X"07",X"34",X"27",X"11",X"83",X"23",X"BB",X"24",X"08",X"10",X"8E",
		X"DF",X"07",X"A6",X"A6",X"A7",X"61",X"1A",X"FF",X"7F",X"C9",X"00",X"34",X"10",X"3A",X"35",X"06",
		X"46",X"56",X"1F",X"98",X"E6",X"64",X"1F",X"02",X"A6",X"61",X"27",X"31",X"24",X"12",X"A8",X"A4",
		X"84",X"0F",X"A8",X"A4",X"A7",X"A4",X"84",X"0F",X"31",X"A9",X"01",X"00",X"6A",X"62",X"27",X"1D",
		X"C6",X"11",X"3D",X"A6",X"62",X"4A",X"27",X"0B",X"E7",X"A4",X"31",X"A9",X"01",X"00",X"4A",X"26",
		X"F4",X"20",X"0A",X"C4",X"F0",X"E8",X"A4",X"C4",X"F0",X"E8",X"A4",X"E7",X"A4",X"86",X"01",X"B7",
		X"C9",X"00",X"35",X"27",X"7E",X"DE",X"52",X"00",X"01",X"08",X"0B",X"0D",X"0F",X"06",X"07",X"AE",
		X"57",X"A6",X"06",X"2B",X"15",X"AE",X"59",X"A6",X"06",X"2B",X"0F",X"AE",X"55",X"A6",X"06",X"2B",
		X"09",X"AE",X"53",X"2A",X"04",X"A6",X"06",X"2B",X"01",X"39",X"10",X"AE",X"06",X"6F",X"06",X"A6",
		X"39",X"85",X"F0",X"26",X"06",X"81",X"0E",X"10",X"26",X"00",X"83",X"81",X"C0",X"10",X"26",X"00",
		X"98",X"10",X"AE",X"2A",X"A6",X"33",X"10",X"2B",X"00",X"96",X"11",X"83",X"9A",X"21",X"10",X"27",
		X"00",X"81",X"A6",X"53",X"2B",X"7D",X"34",X"21",X"1A",X"50",X"10",X"AE",X"A8",X"27",X"10",X"AF",
		X"53",X"EF",X"2A",X"6F",X"25",X"AE",X"55",X"A6",X"03",X"A7",X"23",X"34",X"40",X"EE",X"08",X"EC",
		X"47",X"E3",X"15",X"ED",X"35",X"A6",X"49",X"AB",X"17",X"A7",X"37",X"35",X"40",X"EC",X"51",X"8A",
		X"C0",X"CA",X"03",X"ED",X"51",X"BD",X"5D",X"B9",X"24",X"05",X"CC",X"5D",X"B6",X"ED",X"4A",X"11",
		X"A3",X"61",X"10",X"AE",X"61",X"27",X"23",X"AE",X"C8",X"37",X"EC",X"A8",X"37",X"AF",X"A8",X"37",
		X"ED",X"C8",X"37",X"AE",X"C8",X"27",X"AF",X"A8",X"27",X"6F",X"C8",X"27",X"10",X"AF",X"0A",X"10",
		X"AE",X"53",X"A6",X"0C",X"E6",X"2C",X"A7",X"2C",X"E7",X"0C",X"8D",X"05",X"35",X"21",X"1C",X"FE",
		X"39",X"34",X"20",X"10",X"AE",X"C8",X"37",X"2A",X"05",X"CC",X"D6",X"C5",X"ED",X"22",X"6F",X"C8",
		X"37",X"35",X"A0",X"10",X"AE",X"A8",X"27",X"20",X"0A",X"85",X"80",X"27",X"06",X"10",X"AE",X"2A",
		X"10",X"AE",X"35",X"AE",X"55",X"A6",X"14",X"A0",X"34",X"A7",X"E2",X"A6",X"13",X"A0",X"33",X"AB",
		X"E4",X"47",X"2D",X"04",X"44",X"44",X"20",X"04",X"40",X"44",X"44",X"40",X"A7",X"E4",X"A6",X"11",
		X"A0",X"31",X"34",X"02",X"AE",X"1A",X"A6",X"1B",X"AE",X"3A",X"A0",X"1B",X"47",X"5F",X"AB",X"E0",
		X"2D",X"05",X"44",X"44",X"44",X"20",X"05",X"40",X"44",X"44",X"44",X"40",X"2D",X"06",X"27",X"02",
		X"CB",X"06",X"CB",X"06",X"A6",X"E0",X"2D",X"06",X"27",X"02",X"CB",X"02",X"CB",X"02",X"8E",X"E0",
		X"3E",X"EC",X"85",X"ED",X"47",X"8E",X"E6",X"78",X"BD",X"E6",X"AA",X"1A",X"01",X"39",X"E0",X"9E",
		X"E0",X"50",X"E0",X"6A",X"E0",X"EC",X"00",X"00",X"E1",X"06",X"E0",X"B8",X"E0",X"D2",X"E0",X"84",
		X"05",X"06",X"02",X"02",X"05",X"01",X"01",X"06",X"02",X"05",X"01",X"06",X"02",X"05",X"01",X"06",
		X"02",X"05",X"01",X"06",X"05",X"06",X"05",X"06",X"05",X"00",X"06",X"05",X"06",X"0A",X"0A",X"0A",
		X"06",X"05",X"05",X"05",X"06",X"0A",X"0A",X"06",X"05",X"05",X"06",X"0A",X"02",X"04",X"02",X"04",
		X"02",X"04",X"06",X"00",X"0A",X"09",X"0A",X"06",X"06",X"06",X"0A",X"09",X"09",X"09",X"0A",X"06",
		X"06",X"0A",X"09",X"09",X"0A",X"06",X"02",X"08",X"02",X"08",X"02",X"08",X"0A",X"00",X"05",X"06",
		X"05",X"09",X"09",X"09",X"05",X"06",X"06",X"06",X"05",X"09",X"09",X"05",X"06",X"06",X"05",X"09",
		X"01",X"04",X"01",X"04",X"01",X"04",X"05",X"00",X"09",X"0A",X"09",X"05",X"05",X"05",X"09",X"0A",
		X"0A",X"0A",X"09",X"05",X"05",X"09",X"0A",X"0A",X"09",X"05",X"01",X"08",X"01",X"08",X"01",X"08",
		X"09",X"00",X"0A",X"0A",X"02",X"02",X"09",X"01",X"01",X"0A",X"02",X"09",X"01",X"0A",X"02",X"09",
		X"01",X"0A",X"02",X"09",X"01",X"0A",X"09",X"0A",X"09",X"0A",X"09",X"00",X"01",X"05",X"04",X"04",
		X"09",X"08",X"08",X"05",X"04",X"09",X"08",X"05",X"04",X"09",X"08",X"05",X"04",X"09",X"08",X"05",
		X"09",X"05",X"09",X"05",X"09",X"00",X"02",X"06",X"04",X"04",X"0A",X"08",X"08",X"06",X"04",X"0A",
		X"08",X"06",X"04",X"0A",X"08",X"06",X"04",X"0A",X"08",X"06",X"0A",X"06",X"0A",X"06",X"0A",X"00",
		X"34",X"01",X"1A",X"F0",X"E6",X"25",X"2B",X"78",X"AB",X"22",X"20",X"17",X"34",X"01",X"1A",X"F0",
		X"E6",X"25",X"2B",X"6C",X"1F",X"89",X"84",X"F0",X"C4",X"0F",X"AB",X"23",X"19",X"A7",X"23",X"1F",
		X"98",X"A9",X"22",X"19",X"A7",X"22",X"6C",X"24",X"A6",X"21",X"89",X"00",X"19",X"A7",X"21",X"A6",
		X"A4",X"89",X"00",X"19",X"24",X"02",X"8B",X"10",X"A7",X"A4",X"DC",X"B8",X"27",X"42",X"EC",X"21",
		X"AB",X"26",X"19",X"10",X"A3",X"27",X"25",X"38",X"A6",X"28",X"9B",X"B9",X"19",X"A7",X"28",X"A6",
		X"27",X"99",X"B8",X"19",X"A7",X"27",X"81",X"30",X"25",X"0C",X"8B",X"80",X"19",X"A7",X"27",X"A6",
		X"26",X"8B",X"80",X"19",X"A7",X"26",X"A6",X"25",X"8B",X"01",X"19",X"2B",X"02",X"A7",X"25",X"34",
		X"30",X"8E",X"E6",X"9E",X"BD",X"E6",X"AA",X"C6",X"05",X"BD",X"37",X"B9",X"35",X"30",X"20",X"BE",
		X"35",X"81",X"99",X"10",X"1A",X"22",X"99",X"0C",X"22",X"15",X"E2",X"E8",X"99",X"0D",X"24",X"15",
		X"E2",X"E4",X"99",X"0D",X"26",X"15",X"E2",X"E8",X"99",X"0E",X"28",X"15",X"E2",X"E4",X"99",X"0E",
		X"2A",X"15",X"E2",X"E8",X"99",X"0F",X"2C",X"15",X"E2",X"E4",X"99",X"11",X"34",X"13",X"E2",X"99",
		X"99",X"11",X"37",X"13",X"E2",X"A8",X"00",X"00",X"FF",X"99",X"0F",X"2E",X"15",X"E2",X"E8",X"99",
		X"11",X"34",X"13",X"E2",X"99",X"99",X"11",X"37",X"13",X"E2",X"A8",X"00",X"00",X"FF",X"99",X"19",
		X"1A",X"22",X"99",X"15",X"62",X"15",X"E2",X"E8",X"99",X"16",X"64",X"15",X"E2",X"E4",X"99",X"16",
		X"66",X"15",X"E2",X"E8",X"99",X"17",X"68",X"15",X"E2",X"E4",X"99",X"17",X"6A",X"15",X"E2",X"E8",
		X"99",X"18",X"6C",X"15",X"E2",X"E4",X"99",X"1A",X"5A",X"13",X"E2",X"99",X"99",X"1A",X"5D",X"13",
		X"E2",X"A8",X"00",X"00",X"FF",X"99",X"18",X"6E",X"15",X"E2",X"E8",X"99",X"1A",X"5A",X"13",X"E2",
		X"99",X"99",X"1A",X"5D",X"13",X"E2",X"A8",X"00",X"00",X"FF",X"8E",X"E1",X"A2",X"AF",X"47",X"20",
		X"05",X"8E",X"E1",X"EE",X"AF",X"47",X"30",X"88",X"37",X"AF",X"49",X"10",X"AE",X"47",X"EE",X"22",
		X"10",X"AE",X"02",X"2B",X"0B",X"E6",X"94",X"6E",X"98",X"04",X"AE",X"49",X"30",X"06",X"20",X"E9",
		X"1C",X"AF",X"86",X"04",X"BD",X"D6",X"BA",X"1A",X"50",X"AE",X"47",X"E6",X"94",X"27",X"F1",X"6F",
		X"94",X"1C",X"AF",X"30",X"04",X"E6",X"94",X"26",X"D0",X"30",X"06",X"E6",X"94",X"27",X"08",X"C4",
		X"F0",X"26",X"C6",X"30",X"06",X"20",X"C2",X"30",X"0C",X"E6",X"94",X"27",X"08",X"C4",X"F0",X"26",
		X"B8",X"30",X"06",X"20",X"B4",X"30",X"0C",X"20",X"B0",X"54",X"54",X"54",X"54",X"C1",X"09",X"2E",
		X"03",X"5D",X"26",X"0B",X"C6",X"0A",X"20",X"07",X"C4",X"0F",X"C1",X"09",X"2F",X"01",X"5F",X"86",
		X"17",X"3D",X"34",X"01",X"1A",X"F0",X"E3",X"9F",X"46",X"38",X"C3",X"00",X"02",X"FD",X"CA",X"02",
		X"CC",X"03",X"07",X"FD",X"CA",X"06",X"10",X"BF",X"CA",X"04",X"7F",X"CA",X"01",X"86",X"12",X"B7",
		X"CA",X"00",X"1F",X"30",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"35",X"01",X"86",X"04",X"8E",X"E2",
		X"5A",X"7E",X"D6",X"BC",X"56",X"56",X"56",X"56",X"C4",X"0F",X"C1",X"09",X"22",X"2E",X"86",X"0C",
		X"3D",X"34",X"01",X"1A",X"F0",X"E3",X"9F",X"46",X"40",X"C3",X"00",X"02",X"FD",X"CA",X"02",X"CC",
		X"02",X"05",X"FD",X"CA",X"06",X"10",X"BF",X"CA",X"04",X"7F",X"CA",X"01",X"86",X"12",X"B7",X"CA",
		X"00",X"CC",X"1A",X"44",X"F7",X"CA",X"01",X"B7",X"CA",X"00",X"35",X"01",X"86",X"04",X"8E",X"E2",
		X"5A",X"7E",X"D6",X"BC",X"34",X"01",X"1A",X"F0",X"30",X"02",X"BF",X"CA",X"04",X"BF",X"CA",X"02",
		X"CC",X"0C",X"05",X"FD",X"CA",X"06",X"7F",X"CA",X"01",X"86",X"12",X"B7",X"CA",X"00",X"35",X"81",
		X"0C",X"22",X"CC",X"FF",X"37",X"B7",X"C8",X"0E",X"F7",X"C8",X"0E",X"96",X"39",X"85",X"40",X"26",
		X"01",X"39",X"34",X"01",X"1A",X"50",X"8E",X"3B",X"EB",X"BF",X"CA",X"04",X"BF",X"CA",X"02",X"CC",
		X"15",X"06",X"FD",X"CA",X"06",X"7F",X"C9",X"00",X"E6",X"84",X"F7",X"CA",X"01",X"CC",X"13",X"01",
		X"F7",X"C9",X"00",X"B7",X"CA",X"00",X"8E",X"3C",X"EC",X"CC",X"50",X"44",X"BD",X"46",X"2C",X"B6",
		X"BF",X"32",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"BD",X"46",X"2F",X"35",X"81",X"34",X"12",X"A6",
		X"49",X"27",X"02",X"6A",X"49",X"A6",X"5F",X"10",X"27",X"00",X"CC",X"2A",X"5D",X"6A",X"41",X"26",
		X"4B",X"85",X"40",X"27",X"11",X"84",X"BF",X"A7",X"5F",X"A6",X"E4",X"84",X"C0",X"C4",X"03",X"ED",
		X"61",X"86",X"01",X"7E",X"E4",X"A0",X"A6",X"E4",X"84",X"C0",X"C4",X"03",X"ED",X"61",X"A6",X"5F",
		X"84",X"7F",X"A7",X"5F",X"64",X"61",X"64",X"61",X"64",X"61",X"64",X"61",X"E6",X"62",X"EA",X"61",
		X"27",X"0F",X"10",X"8E",X"E4",X"D8",X"44",X"24",X"04",X"10",X"8E",X"E4",X"E8",X"E6",X"A5",X"E7",
		X"42",X"A6",X"42",X"27",X"48",X"86",X"02",X"A7",X"41",X"32",X"63",X"39",X"85",X"40",X"27",X"F9",
		X"EA",X"E4",X"C5",X"C3",X"26",X"F3",X"6F",X"5F",X"20",X"EF",X"6A",X"41",X"26",X"2C",X"34",X"01",
		X"1A",X"50",X"A6",X"5F",X"44",X"24",X"07",X"AE",X"59",X"10",X"AE",X"5D",X"20",X"05",X"AE",X"57",
		X"10",X"AE",X"5B",X"2A",X"4E",X"6C",X"25",X"BD",X"D8",X"D8",X"35",X"01",X"8E",X"E6",X"72",X"BD",
		X"E6",X"AA",X"E6",X"25",X"E1",X"42",X"24",X"05",X"6C",X"41",X"32",X"63",X"39",X"A6",X"5F",X"44",
		X"25",X"11",X"AE",X"57",X"10",X"AE",X"5B",X"2A",X"24",X"4F",X"5F",X"ED",X"5B",X"1F",X"20",X"84",
		X"7F",X"20",X"0D",X"AE",X"59",X"10",X"AE",X"5D",X"2A",X"13",X"4F",X"5F",X"ED",X"5D",X"1F",X"20",
		X"6D",X"C8",X"2F",X"27",X"05",X"ED",X"C8",X"31",X"20",X"03",X"ED",X"C8",X"2F",X"6F",X"02",X"6F",
		X"5F",X"20",X"66",X"35",X"01",X"20",X"F6",X"A6",X"E4",X"84",X"C0",X"26",X"04",X"C4",X"03",X"27",
		X"58",X"C4",X"03",X"ED",X"61",X"CC",X"02",X"81",X"10",X"AE",X"5D",X"2B",X"06",X"10",X"AE",X"5B",
		X"2A",X"47",X"5C",X"E7",X"5F",X"E6",X"39",X"54",X"C1",X"05",X"26",X"10",X"10",X"AE",X"5B",X"2A",
		X"3B",X"E6",X"39",X"54",X"C1",X"05",X"27",X"34",X"C6",X"82",X"E7",X"5F",X"C6",X"14",X"E7",X"49",
		X"A7",X"41",X"64",X"61",X"64",X"61",X"64",X"61",X"64",X"61",X"A6",X"62",X"AA",X"61",X"10",X"8E",
		X"E4",X"D8",X"AE",X"57",X"E6",X"5F",X"C5",X"01",X"27",X"06",X"10",X"8E",X"E4",X"E8",X"AE",X"59",
		X"A6",X"A6",X"A7",X"42",X"6C",X"02",X"BD",X"DC",X"73",X"32",X"63",X"39",X"AB",X"49",X"A7",X"41",
		X"E6",X"5F",X"CA",X"40",X"E7",X"5F",X"20",X"F1",X"00",X"06",X"02",X"00",X"00",X"07",X"01",X"00",
		X"04",X"05",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"00",X"00",X"01",X"07",X"00",
		X"04",X"03",X"05",X"00",X"00",X"00",X"00",X"00",X"E5",X"06",X"E5",X"06",X"E5",X"06",X"E5",X"26",
		X"E5",X"26",X"E5",X"06",X"E5",X"26",X"00",X"00",X"FC",X"88",X"01",X"39",X"FD",X"8D",X"01",X"6C",
		X"00",X"00",X"01",X"39",X"02",X"73",X"00",X"00",X"03",X"78",X"FE",X"C7",X"02",X"73",X"FE",X"94",
		X"00",X"00",X"FE",X"C7",X"FD",X"8D",X"00",X"00",X"FC",X"E8",X"01",X"17",X"FD",X"D1",X"01",X"8C",
		X"00",X"00",X"01",X"17",X"02",X"2F",X"00",X"00",X"03",X"18",X"FE",X"E9",X"02",X"2F",X"FE",X"74",
		X"00",X"00",X"FE",X"E9",X"FD",X"D1",X"86",X"C8",X"BD",X"D6",X"BA",X"CC",X"A1",X"20",X"8D",X"6C",
		X"26",X"F4",X"8D",X"68",X"27",X"FC",X"86",X"0F",X"BD",X"D6",X"BA",X"CC",X"20",X"68",X"8D",X"5C",
		X"26",X"E4",X"8D",X"58",X"27",X"FC",X"86",X"0F",X"BD",X"D6",X"BA",X"CC",X"41",X"82",X"8D",X"4C",
		X"26",X"D4",X"1A",X"50",X"CC",X"00",X"FF",X"FD",X"C0",X"00",X"BD",X"DD",X"0F",X"CE",X"E5",X"D6",
		X"8E",X"10",X"30",X"34",X"10",X"C6",X"11",X"A6",X"C0",X"88",X"9B",X"80",X"35",X"2B",X"10",X"27",
		X"05",X"BD",X"46",X"20",X"20",X"F1",X"AE",X"E4",X"30",X"88",X"10",X"AF",X"E4",X"20",X"E8",X"8E",
		X"1B",X"E6",X"86",X"39",X"B7",X"CB",X"FF",X"BD",X"E6",X"42",X"84",X"41",X"C4",X"82",X"10",X"83",
		X"41",X"82",X"27",X"EB",X"30",X"1F",X"26",X"EA",X"6E",X"9F",X"FF",X"FE",X"ED",X"47",X"35",X"06",
		X"ED",X"49",X"86",X"08",X"BD",X"D6",X"BA",X"8D",X"79",X"A4",X"47",X"E4",X"48",X"1F",X"01",X"EC",
		X"47",X"AC",X"47",X"6E",X"D8",X"09",X"C8",X"DC",X"D3",X"C9",X"A4",X"D3",X"C9",X"A4",X"C9",X"D4",
		X"D0",X"DB",X"C8",X"F8",X"AE",X"D8",X"DF",X"C9",X"D3",X"DD",X"D6",X"DF",X"D8",X"A4",X"DA",X"C3",
		X"A4",X"CD",X"D3",X"D0",X"D0",X"D3",X"DB",X"D7",X"C9",X"A4",X"DF",X"D0",X"DF",X"D9",X"C8",X"CA",
		X"D5",X"D6",X"D3",X"D9",X"C9",X"A4",X"D3",X"D6",X"D9",X"F8",X"AE",X"C4",X"D9",X"FB",X"A4",X"AD",
		X"A5",X"A6",X"AC",X"A4",X"CD",X"D3",X"D0",X"D0",X"D3",X"DB",X"D7",X"C9",X"A4",X"DF",X"D0",X"DF",
		X"D9",X"C8",X"CA",X"D5",X"D6",X"D3",X"D9",X"C9",X"A4",X"D3",X"D6",X"D9",X"F8",X"AE",X"DB",X"D0",
		X"D0",X"A4",X"CA",X"D3",X"DD",X"DC",X"C8",X"C9",X"A4",X"CA",X"DF",X"C9",X"DF",X"CA",X"CE",X"DF",
		X"D8",X"2E",X"34",X"01",X"1A",X"50",X"86",X"08",X"BA",X"C8",X"07",X"B7",X"C8",X"07",X"B6",X"C8",
		X"04",X"C6",X"F7",X"F4",X"C8",X"07",X"F7",X"C8",X"07",X"F6",X"C8",X"04",X"35",X"81",X"0A",X"75",
		X"0F",X"0A",X"74",X"0F",X"14",X"73",X"0F",X"1E",X"71",X"0F",X"28",X"78",X"14",X"28",X"E4",X"05",
		X"64",X"0F",X"28",X"61",X"0C",X"32",X"70",X"0F",X"32",X"76",X"0F",X"3C",X"60",X"0C",X"46",X"6F",
		X"23",X"46",X"F8",X"19",X"72",X"05",X"46",X"72",X"05",X"50",X"73",X"0F",X"5A",X"EB",X"F0",X"3F",
		X"B4",X"5B",X"E4",X"01",X"64",X"0F",X"64",X"72",X"04",X"6E",X"F7",X"15",X"6E",X"1E",X"78",X"77",
		X"28",X"C8",X"7B",X"01",X"D2",X"68",X"80",X"DC",X"72",X"08",X"34",X"07",X"1A",X"F0",X"A6",X"80",
		X"2B",X"07",X"D6",X"39",X"53",X"C5",X"03",X"27",X"10",X"D6",X"64",X"27",X"04",X"91",X"65",X"25",
		X"08",X"97",X"65",X"86",X"01",X"97",X"64",X"9F",X"66",X"35",X"87",X"27",X"2B",X"1B",X"66",X"2A",
		X"2B",X"1B",X"AB",X"33",X"2B",X"1B",X"AB",X"58",X"2B",X"1B",X"EC",X"61",X"2B",X"1B",X"EC",X"6A",
		X"2B",X"1C",X"AA",X"27",X"2B",X"1B",X"7D",X"2A",X"2B",X"1B",X"EC",X"33",X"2B",X"1B",X"EC",X"58",
		X"2B",X"1B",X"AB",X"61",X"2B",X"1B",X"AB",X"6A",X"2B",X"1C",X"8C",X"27",X"2B",X"1B",X"94",X"2A",
		X"2B",X"1C",X"2D",X"33",X"2B",X"1C",X"2D",X"58",X"2B",X"1C",X"2D",X"61",X"2B",X"1C",X"2D",X"6A",
		X"2B",X"1C",X"6E",X"CC",X"D0",X"0D",X"B7",X"3C",X"33",X"F7",X"57",X"33",X"8E",X"00",X"78",X"10",
		X"8E",X"00",X"09",X"CE",X"17",X"E2",X"BD",X"DE",X"4E",X"8E",X"E6",X"5E",X"BD",X"E6",X"AA",X"8E",
		X"E7",X"E9",X"10",X"AE",X"81",X"BD",X"E7",X"62",X"8C",X"E7",X"F3",X"25",X"F5",X"86",X"0F",X"BD",
		X"D6",X"BA",X"96",X"68",X"27",X"F7",X"8E",X"E6",X"61",X"BD",X"E6",X"AA",X"8E",X"E7",X"F3",X"10",
		X"AE",X"81",X"BD",X"E7",X"62",X"8C",X"E7",X"FD",X"25",X"F5",X"86",X"0F",X"8E",X"E7",X"29",X"7E",
		X"D6",X"BC",X"34",X"01",X"1A",X"50",X"EC",X"A1",X"FD",X"CA",X"06",X"EC",X"A4",X"FD",X"CA",X"04",
		X"31",X"23",X"10",X"BF",X"CA",X"02",X"A6",X"3F",X"B7",X"CA",X"00",X"35",X"81",X"AE",X"C1",X"10",
		X"AE",X"C1",X"1A",X"50",X"EC",X"A4",X"FD",X"CA",X"06",X"31",X"22",X"10",X"BF",X"CA",X"02",X"BF",
		X"CA",X"04",X"86",X"02",X"B7",X"CA",X"00",X"1C",X"AF",X"39",X"CE",X"E6",X"CB",X"8D",X"DE",X"11",
		X"83",X"E6",X"E3",X"26",X"F8",X"86",X"03",X"BD",X"D6",X"BA",X"CE",X"E6",X"E3",X"8D",X"CE",X"11",
		X"83",X"E6",X"FB",X"26",X"F8",X"86",X"03",X"BD",X"D6",X"BA",X"CE",X"E6",X"FB",X"8D",X"BE",X"11",
		X"83",X"E7",X"13",X"26",X"F8",X"86",X"03",X"BD",X"D6",X"BA",X"96",X"68",X"26",X"CC",X"A6",X"47",
		X"26",X"06",X"6C",X"47",X"86",X"10",X"A7",X"48",X"6A",X"48",X"26",X"BE",X"86",X"06",X"BD",X"D6",
		X"BA",X"96",X"68",X"27",X"F7",X"6F",X"47",X"20",X"B1",X"1A",X"95",X"1A",X"CF",X"1A",X"F7",X"1B",
		X"27",X"1B",X"59",X"1A",X"78",X"1A",X"B2",X"1A",X"EC",X"1B",X"02",X"1B",X"4C",X"34",X"76",X"CC",
		X"6E",X"11",X"CE",X"40",X"60",X"BD",X"E8",X"8D",X"A6",X"E4",X"4C",X"BD",X"D9",X"17",X"85",X"F0",
		X"26",X"02",X"8A",X"F0",X"CE",X"4F",X"60",X"BD",X"E8",X"83",X"E6",X"E4",X"C1",X"04",X"24",X"1B",
		X"BD",X"D6",X"8B",X"E9",X"10",X"38",X"86",X"CD",X"10",X"8E",X"21",X"A0",X"C1",X"03",X"26",X"06",
		X"86",X"69",X"10",X"8E",X"2D",X"80",X"A7",X"08",X"10",X"AF",X"09",X"C0",X"06",X"24",X"FC",X"CB",
		X"06",X"86",X"09",X"3D",X"10",X"8E",X"E8",X"A0",X"31",X"A5",X"C1",X"12",X"27",X"0A",X"EC",X"A4",
		X"6D",X"E4",X"26",X"16",X"C6",X"00",X"20",X"12",X"96",X"CA",X"CE",X"E8",X"D6",X"33",X"C6",X"8B",
		X"04",X"81",X"10",X"25",X"01",X"4F",X"97",X"CA",X"EC",X"C4",X"D7",X"73",X"C6",X"11",X"EE",X"22",
		X"8D",X"1B",X"A6",X"26",X"27",X"06",X"C6",X"22",X"EE",X"27",X"8D",X"11",X"AE",X"24",X"BD",X"E6",
		X"AA",X"35",X"F6",X"97",X"3D",X"BD",X"D6",X"8B",X"E8",X"EB",X"00",X"20",X"08",X"97",X"3D",X"BD",
		X"D6",X"8B",X"E8",X"E6",X"35",X"96",X"3D",X"ED",X"07",X"EF",X"09",X"86",X"1E",X"A7",X"0B",X"39",
		X"60",X"80",X"3C",X"70",X"E6",X"A1",X"00",X"21",X"80",X"62",X"03",X"3B",X"70",X"E6",X"A1",X"66",
		X"30",X"80",X"61",X"04",X"38",X"70",X"E6",X"A1",X"6A",X"2E",X"80",X"D6",X"05",X"33",X"70",X"E6",
		X"A1",X"00",X"2D",X"80",X"D5",X"80",X"3D",X"70",X"E6",X"A1",X"00",X"45",X"70",X"D4",X"00",X"3A",
		X"70",X"E6",X"A1",X"D3",X"32",X"80",X"61",X"04",X"38",X"70",X"63",X"02",X"3B",X"70",X"65",X"01",
		X"37",X"70",X"64",X"00",X"36",X"70",X"CC",X"46",X"23",X"20",X"08",X"CC",X"46",X"26",X"20",X"03",
		X"CC",X"46",X"2C",X"ED",X"4D",X"86",X"03",X"BD",X"D6",X"BA",X"EC",X"47",X"AE",X"49",X"AD",X"D8",
		X"0D",X"6A",X"4B",X"26",X"F0",X"A6",X"47",X"5F",X"AE",X"49",X"AD",X"D8",X"0D",X"7E",X"D6",X"C5",
		X"86",X"0F",X"A7",X"47",X"6A",X"47",X"10",X"27",X"ED",X"AB",X"BD",X"D6",X"8B",X"E8",X"E6",X"27",
		X"A6",X"48",X"C6",X"22",X"ED",X"07",X"EC",X"49",X"ED",X"09",X"86",X"04",X"A7",X"0B",X"86",X"0F",
		X"8E",X"E9",X"14",X"7E",X"D6",X"BC",X"2D",X"3B",X"03",X"B0",X"2D",X"3B",X"03",X"45",X"2F",X"2D",
		X"90",X"45",X"2F",X"2D",X"90",X"B0",X"31",X"1F",X"42",X"33",X"2D",X"D5",X"03",X"B0",X"2D",X"D5",
		X"03",X"45",X"2F",X"C7",X"8B",X"45",X"2F",X"C7",X"8B",X"B0",X"31",X"51",X"42",X"33",X"2D",X"D5",
		X"03",X"B0",X"2D",X"D5",X"03",X"45",X"2F",X"C7",X"8B",X"45",X"2F",X"C7",X"8B",X"B0",X"31",X"C3",
		X"42",X"33",X"34",X"15",X"8E",X"98",X"9E",X"E6",X"86",X"26",X"06",X"C6",X"1E",X"E7",X"86",X"35",
		X"95",X"C1",X"19",X"24",X"FA",X"C6",X"19",X"20",X"F4",X"4F",X"5F",X"ED",X"47",X"ED",X"49",X"A7",
		X"4B",X"4F",X"33",X"47",X"8E",X"98",X"9E",X"E6",X"86",X"27",X"2E",X"6A",X"86",X"26",X"07",X"C6",
		X"80",X"E7",X"C6",X"5F",X"20",X"1E",X"C1",X"05",X"25",X"12",X"C1",X"19",X"24",X"0E",X"C6",X"02",
		X"6D",X"C6",X"2B",X"10",X"C6",X"80",X"E7",X"C6",X"C6",X"02",X"20",X"08",X"C6",X"01",X"6D",X"C6",
		X"2A",X"02",X"6F",X"C6",X"8E",X"98",X"AD",X"E7",X"86",X"4C",X"81",X"05",X"26",X"C6",X"86",X"03",
		X"8E",X"E9",X"91",X"7E",X"D6",X"BC",X"86",X"F0",X"BD",X"D6",X"BA",X"86",X"1E",X"BD",X"D6",X"BA",
		X"86",X"01",X"BD",X"D6",X"BA",X"D6",X"86",X"27",X"F2",X"96",X"39",X"43",X"85",X"03",X"27",X"E6",
		X"44",X"24",X"07",X"BE",X"99",X"86",X"E6",X"11",X"26",X"0A",X"44",X"24",X"E3",X"BE",X"99",X"CE",
		X"E6",X"11",X"27",X"D7",X"BD",X"EA",X"F2",X"2B",X"D2",X"10",X"AF",X"4B",X"8E",X"98",X"A3",X"6C",
		X"86",X"BD",X"E9",X"72",X"86",X"1E",X"BD",X"D6",X"BA",X"AE",X"4B",X"A6",X"16",X"10",X"8E",X"98",
		X"A3",X"6A",X"A6",X"A6",X"15",X"E6",X"17",X"34",X"06",X"CE",X"9A",X"21",X"6F",X"C8",X"22",X"63",
		X"C8",X"26",X"CC",X"FF",X"FF",X"ED",X"51",X"86",X"01",X"A7",X"C8",X"19",X"FC",X"99",X"86",X"ED",
		X"C8",X"17",X"6F",X"C8",X"1A",X"6F",X"C8",X"1B",X"CC",X"EB",X"B3",X"ED",X"4A",X"86",X"FF",X"A7",
		X"C8",X"23",X"6F",X"C8",X"24",X"6F",X"C8",X"10",X"1A",X"50",X"EC",X"E4",X"BD",X"73",X"75",X"FE",
		X"9A",X"1A",X"8E",X"9A",X"1E",X"BD",X"EF",X"4A",X"FE",X"9A",X"18",X"8E",X"9A",X"1C",X"BD",X"EF",
		X"4A",X"1C",X"AF",X"32",X"62",X"86",X"01",X"BD",X"D6",X"BA",X"CE",X"9A",X"21",X"AE",X"55",X"A6",
		X"11",X"27",X"11",X"0A",X"BB",X"26",X"0D",X"B6",X"99",X"07",X"97",X"BB",X"BD",X"D6",X"8B",X"69",
		X"87",X"33",X"AE",X"55",X"BD",X"6F",X"67",X"A6",X"C8",X"23",X"2B",X"0A",X"A6",X"C8",X"24",X"2B",
		X"27",X"BD",X"71",X"A3",X"20",X"CF",X"BD",X"74",X"6E",X"AE",X"47",X"27",X"0D",X"84",X"F0",X"AA",
		X"80",X"6D",X"84",X"26",X"03",X"8E",X"00",X"00",X"AF",X"47",X"AE",X"55",X"A4",X"51",X"E4",X"52",
		X"BD",X"70",X"22",X"BD",X"E3",X"8D",X"20",X"AD",X"1A",X"F0",X"AE",X"5D",X"8D",X"0F",X"AF",X"5D",
		X"AE",X"5B",X"8D",X"09",X"AF",X"5B",X"1C",X"AF",X"6F",X"5F",X"7E",X"E9",X"E0",X"2A",X"03",X"BD",
		X"D7",X"84",X"8E",X"00",X"00",X"39",X"0F",X"00",X"BF",X"0F",X"01",X"54",X"80",X"02",X"54",X"80",
		X"03",X"BF",X"34",X"15",X"1A",X"F0",X"0F",X"92",X"20",X"0E",X"34",X"15",X"1A",X"F0",X"0F",X"92",
		X"96",X"A7",X"97",X"97",X"26",X"02",X"0C",X"92",X"DC",X"A3",X"DD",X"93",X"4D",X"26",X"02",X"0C",
		X"92",X"5D",X"26",X"02",X"0C",X"92",X"DC",X"A5",X"DD",X"95",X"4D",X"26",X"02",X"0C",X"92",X"5D",
		X"26",X"02",X"0C",X"92",X"BE",X"99",X"86",X"8D",X"44",X"BE",X"99",X"CE",X"8D",X"3F",X"BE",X"9A",
		X"16",X"8D",X"3A",X"9E",X"77",X"2A",X"02",X"8D",X"38",X"9E",X"79",X"2A",X"02",X"8D",X"32",X"BD",
		X"5D",X"BF",X"D6",X"92",X"27",X"1D",X"3D",X"C6",X"FF",X"8E",X"98",X"93",X"5C",X"6D",X"85",X"26",
		X"FB",X"4A",X"2A",X"F8",X"1F",X"98",X"34",X"04",X"58",X"EB",X"E0",X"10",X"8E",X"EA",X"F1",X"31",
		X"A5",X"20",X"06",X"10",X"8E",X"00",X"00",X"86",X"FF",X"35",X"15",X"4D",X"39",X"AC",X"55",X"27",
		X"1E",X"E6",X"11",X"27",X"1A",X"A6",X"13",X"81",X"79",X"23",X"1E",X"81",X"97",X"25",X"10",X"C1",
		X"2D",X"23",X"0D",X"C1",X"63",X"25",X"08",X"96",X"96",X"26",X"04",X"0C",X"96",X"0A",X"92",X"39",
		X"96",X"93",X"26",X"FB",X"0C",X"93",X"0A",X"92",X"39",X"C1",X"2D",X"23",X"0D",X"C1",X"63",X"25",
		X"EE",X"96",X"95",X"26",X"EA",X"0C",X"95",X"0A",X"92",X"39",X"96",X"94",X"26",X"E1",X"0C",X"94",
		X"0A",X"92",X"39",X"D6",X"86",X"27",X"22",X"6A",X"C8",X"19",X"26",X"52",X"86",X"0F",X"A7",X"C8",
		X"19",X"96",X"39",X"44",X"25",X"08",X"10",X"BE",X"99",X"86",X"E6",X"31",X"26",X"0E",X"10",X"BE",
		X"99",X"CE",X"E6",X"31",X"27",X"03",X"44",X"24",X"31",X"7E",X"EC",X"5B",X"44",X"25",X"27",X"10",
		X"BE",X"99",X"CE",X"E6",X"31",X"27",X"1F",X"BD",X"ED",X"56",X"34",X"06",X"10",X"BE",X"99",X"86",
		X"BD",X"ED",X"56",X"10",X"A3",X"E4",X"23",X"06",X"EC",X"E4",X"10",X"BE",X"99",X"CE",X"32",X"62",
		X"10",X"AF",X"C8",X"17",X"20",X"0F",X"10",X"BE",X"99",X"86",X"10",X"AF",X"C8",X"17",X"10",X"AE",
		X"C8",X"17",X"BD",X"ED",X"56",X"93",X"E8",X"25",X"0B",X"C6",X"05",X"BD",X"ED",X"78",X"BD",X"EF",
		X"64",X"7E",X"79",X"70",X"6D",X"5B",X"26",X"09",X"6D",X"5D",X"26",X"0A",X"4F",X"5F",X"7E",X"79",
		X"70",X"CC",X"EC",X"43",X"20",X"03",X"CC",X"EC",X"4C",X"ED",X"4A",X"BD",X"78",X"DC",X"ED",X"4C",
		X"7E",X"79",X"70",X"A6",X"5B",X"27",X"09",X"EC",X"4C",X"7E",X"79",X"70",X"A6",X"5D",X"26",X"F7",
		X"CC",X"EB",X"B3",X"ED",X"4A",X"6F",X"C8",X"22",X"7E",X"EB",X"B3",X"86",X"01",X"A7",X"C8",X"19",
		X"6F",X"C8",X"22",X"C6",X"FF",X"E7",X"C8",X"12",X"D6",X"86",X"27",X"18",X"96",X"39",X"44",X"25",
		X"08",X"10",X"BE",X"99",X"86",X"E6",X"31",X"26",X"D7",X"44",X"25",X"08",X"10",X"BE",X"99",X"CE",
		X"E6",X"31",X"26",X"CC",X"CC",X"EC",X"8C",X"ED",X"4A",X"BD",X"EC",X"DB",X"A6",X"C8",X"23",X"2A",
		X"9B",X"6A",X"C8",X"16",X"2F",X"D2",X"A6",X"47",X"27",X"05",X"86",X"FF",X"A7",X"C8",X"12",X"10",
		X"AE",X"C8",X"13",X"5F",X"BD",X"ED",X"78",X"BD",X"EF",X"64",X"34",X"05",X"1A",X"F0",X"4D",X"26",
		X"09",X"E6",X"47",X"26",X"05",X"E6",X"36",X"E7",X"C8",X"23",X"35",X"05",X"7E",X"79",X"70",X"6F",
		X"C8",X"22",X"C6",X"FF",X"E7",X"C8",X"12",X"CC",X"EC",X"CE",X"ED",X"4A",X"8D",X"0D",X"A6",X"53",
		X"10",X"2A",X"87",X"DB",X"6A",X"C8",X"16",X"2F",X"EE",X"20",X"BB",X"C6",X"0F",X"E7",X"C8",X"16",
		X"10",X"8E",X"FF",X"FF",X"34",X"76",X"10",X"8E",X"EA",X"F1",X"A6",X"36",X"8E",X"98",X"A3",X"E6",
		X"86",X"26",X"36",X"AE",X"55",X"8D",X"5F",X"ED",X"E4",X"BE",X"99",X"CE",X"11",X"83",X"99",X"D9",
		X"26",X"03",X"BE",X"9A",X"16",X"8D",X"4F",X"A3",X"E4",X"25",X"1E",X"BE",X"99",X"86",X"11",X"83",
		X"99",X"91",X"26",X"03",X"BE",X"9A",X"16",X"8D",X"3D",X"A3",X"E4",X"25",X"0C",X"EC",X"E4",X"10",
		X"A3",X"64",X"22",X"05",X"ED",X"64",X"10",X"AF",X"66",X"31",X"23",X"10",X"8C",X"EA",X"FA",X"23",
		X"B9",X"35",X"16",X"35",X"26",X"83",X"FF",X"FF",X"27",X"0A",X"86",X"FF",X"A7",X"C8",X"12",X"10",
		X"AF",X"C8",X"13",X"39",X"A6",X"C8",X"12",X"2A",X"0C",X"BD",X"EA",X"F2",X"2B",X"07",X"A7",X"C8",
		X"12",X"10",X"AF",X"C8",X"13",X"39",X"A6",X"11",X"27",X"1A",X"A6",X"35",X"A0",X"15",X"22",X"01",
		X"40",X"1F",X"89",X"3D",X"ED",X"E3",X"E6",X"37",X"E0",X"17",X"22",X"01",X"50",X"54",X"1F",X"98",
		X"3D",X"E3",X"E1",X"39",X"CC",X"FF",X"FF",X"39",X"4F",X"34",X"32",X"EB",X"37",X"C1",X"D5",X"23",
		X"02",X"C6",X"D5",X"34",X"04",X"E6",X"17",X"BC",X"9A",X"16",X"26",X"02",X"CB",X"0A",X"E0",X"E0",
		X"27",X"11",X"22",X"09",X"50",X"54",X"54",X"27",X"0A",X"8A",X"02",X"20",X"06",X"54",X"54",X"27",
		X"02",X"8A",X"01",X"E7",X"C8",X"21",X"E6",X"15",X"E0",X"35",X"27",X"12",X"22",X"0B",X"50",X"54",
		X"27",X"0C",X"8A",X"08",X"20",X"08",X"7E",X"EF",X"44",X"54",X"27",X"02",X"8A",X"04",X"E7",X"C8",
		X"20",X"A7",X"E4",X"27",X"F1",X"10",X"9E",X"7E",X"27",X"EC",X"C6",X"FD",X"A6",X"15",X"8B",X"FE",
		X"A0",X"35",X"22",X"13",X"40",X"81",X"17",X"22",X"DD",X"81",X"13",X"24",X"1A",X"A6",X"15",X"81",
		X"0F",X"27",X"14",X"CB",X"02",X"20",X"10",X"81",X"16",X"22",X"CB",X"5C",X"81",X"12",X"24",X"07",
		X"A6",X"15",X"81",X"80",X"27",X"01",X"5C",X"A6",X"34",X"80",X"13",X"A0",X"17",X"23",X"0E",X"81",
		X"1E",X"22",X"B3",X"CB",X"03",X"81",X"15",X"24",X"11",X"CB",X"06",X"20",X"0D",X"40",X"81",X"1E",
		X"22",X"A4",X"CB",X"06",X"81",X"15",X"24",X"02",X"CB",X"03",X"C1",X"08",X"10",X"26",X"00",X"B0",
		X"86",X"08",X"E6",X"15",X"C0",X"02",X"E1",X"35",X"22",X"01",X"44",X"E6",X"34",X"C0",X"13",X"E1",
		X"17",X"25",X"02",X"8A",X"01",X"7E",X"EF",X"44",X"01",X"02",X"00",X"04",X"08",X"10",X"00",X"20",
		X"40",X"80",X"80",X"10",X"92",X"40",X"08",X"49",X"E0",X"1C",X"FF",X"FF",X"7F",X"FF",X"FF",X"F7",
		X"BF",X"EF",X"FF",X"FF",X"EF",X"FF",X"FF",X"BF",X"7F",X"F7",X"08",X"02",X"08",X"01",X"04",X"04",
		X"01",X"02",X"02",X"04",X"04",X"08",X"01",X"08",X"02",X"01",X"57",X"56",X"73",X"54",X"53",X"70",
		X"3C",X"3B",X"02",X"04",X"04",X"08",X"01",X"08",X"02",X"01",X"02",X"02",X"00",X"01",X"01",X"08",
		X"08",X"00",X"04",X"04",X"86",X"01",X"E6",X"34",X"C0",X"13",X"C1",X"C0",X"24",X"38",X"10",X"AE",
		X"63",X"E1",X"37",X"22",X"31",X"86",X"02",X"20",X"2D",X"C6",X"38",X"A6",X"C8",X"21",X"A1",X"C8",
		X"20",X"22",X"02",X"C6",X"3D",X"A6",X"85",X"81",X"02",X"26",X"1B",X"E6",X"34",X"C0",X"13",X"C1",
		X"C0",X"25",X"13",X"86",X"01",X"20",X"0F",X"86",X"08",X"E6",X"35",X"CB",X"02",X"10",X"AE",X"63",
		X"E1",X"35",X"22",X"02",X"86",X"04",X"A7",X"E4",X"C6",X"30",X"A5",X"85",X"27",X"2E",X"20",X"49",
		X"8E",X"EE",X"37",X"A6",X"E4",X"84",X"0F",X"A6",X"86",X"CB",X"0B",X"A4",X"85",X"27",X"68",X"30",
		X"85",X"E6",X"C8",X"22",X"26",X"40",X"C6",X"08",X"A4",X"85",X"26",X"17",X"C6",X"18",X"A6",X"85",
		X"81",X"02",X"26",X"08",X"A6",X"34",X"80",X"13",X"81",X"C0",X"24",X"1D",X"C6",X"01",X"E7",X"C8",
		X"22",X"20",X"23",X"C6",X"10",X"A4",X"85",X"26",X"17",X"C6",X"20",X"A6",X"85",X"81",X"02",X"26",
		X"08",X"A6",X"34",X"80",X"13",X"81",X"C0",X"24",X"E3",X"C6",X"FF",X"E7",X"C8",X"22",X"20",X"06",
		X"C6",X"28",X"A6",X"85",X"6E",X"86",X"C6",X"18",X"A6",X"C8",X"22",X"2A",X"02",X"C6",X"20",X"A6",
		X"85",X"81",X"02",X"26",X"0B",X"AE",X"61",X"E6",X"17",X"C1",X"D6",X"25",X"03",X"60",X"C8",X"22",
		X"A7",X"E4",X"20",X"03",X"6F",X"C8",X"22",X"5F",X"35",X"B2",X"34",X"50",X"BD",X"D7",X"50",X"9F",
		X"2A",X"86",X"00",X"BD",X"D6",X"45",X"EE",X"62",X"A6",X"59",X"BD",X"D5",X"5A",X"AE",X"F4",X"BD",
		X"D8",X"C6",X"35",X"D0",X"0D",X"E6",X"27",X"1C",X"6D",X"C8",X"26",X"2A",X"06",X"85",X"03",X"26",
		X"11",X"20",X"06",X"85",X"0C",X"26",X"05",X"20",X"06",X"63",X"C8",X"26",X"84",X"FC",X"39",X"63",
		X"C8",X"26",X"84",X"F3",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D7",X"AE",X"D7",X"AE",X"D7",X"AE",X"D7",X"AE",X"D9",X"2E",X"D7",X"AE",X"D7",X"AE",X"D7",X"AE",
		X"7E",X"F0",X"22",X"7E",X"F3",X"3F",X"7E",X"F4",X"6C",X"7E",X"F9",X"5C",X"7E",X"FF",X"23",X"7E",
		X"FF",X"97",X"00",X"F9",X"07",X"28",X"2F",X"00",X"A4",X"15",X"C7",X"FF",X"38",X"17",X"CC",X"81",
		X"81",X"2F",X"1A",X"FF",X"10",X"CE",X"BF",X"00",X"7F",X"C8",X"0D",X"7F",X"C8",X"0C",X"86",X"3C",
		X"B7",X"C8",X"0D",X"7F",X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"3C",X"B7",X"C8",X"0F",
		X"86",X"C0",X"B7",X"C8",X"0E",X"86",X"01",X"B7",X"C9",X"00",X"8E",X"F0",X"12",X"10",X"8E",X"C0",
		X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"F0",X"22",X"25",X"F7",X"86",X"02",X"10",X"8E",X"F0",X"65",
		X"8E",X"00",X"00",X"20",X"3A",X"10",X"8E",X"F0",X"6C",X"7E",X"F2",X"8B",X"86",X"34",X"B7",X"C8",
		X"0D",X"B7",X"C8",X"0F",X"7F",X"C8",X"0E",X"86",X"BF",X"1F",X"8B",X"10",X"CE",X"BF",X"00",X"BD",
		X"37",X"BC",X"86",X"05",X"8E",X"30",X"70",X"C6",X"99",X"BD",X"46",X"23",X"86",X"06",X"8E",X"3A",
		X"90",X"C6",X"99",X"BD",X"46",X"23",X"10",X"8E",X"FF",X"97",X"86",X"07",X"7E",X"F1",X"CB",X"1A",
		X"3F",X"7F",X"C9",X"00",X"1F",X"8B",X"1F",X"10",X"1F",X"03",X"8E",X"00",X"00",X"53",X"C5",X"09",
		X"26",X"05",X"53",X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",
		X"44",X"56",X"ED",X"81",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"B9",
		X"C1",X"FF",X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",X"5F",X"1E",X"10",
		X"8C",X"C0",X"00",X"26",X"C8",X"1F",X"30",X"8E",X"00",X"00",X"53",X"C5",X"09",X"26",X"05",X"53",
		X"46",X"56",X"20",X"0B",X"53",X"C5",X"09",X"26",X"04",X"46",X"56",X"20",X"02",X"44",X"56",X"10",
		X"A3",X"81",X"26",X"43",X"1E",X"10",X"5D",X"26",X"15",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"B9",
		X"C1",X"FF",X"26",X"09",X"F6",X"C8",X"0C",X"C5",X"02",X"27",X"02",X"6E",X"A4",X"5F",X"1E",X"10",
		X"8C",X"C0",X"00",X"26",X"C5",X"1F",X"03",X"1F",X"B8",X"81",X"FF",X"26",X"05",X"1F",X"30",X"7E",
		X"F0",X"AA",X"4A",X"1F",X"8B",X"81",X"80",X"27",X"07",X"4D",X"1F",X"30",X"10",X"26",X"FF",X"6A",
		X"C6",X"01",X"F7",X"C9",X"00",X"6E",X"A4",X"30",X"1E",X"A8",X"84",X"E8",X"01",X"4D",X"26",X"07",
		X"5D",X"26",X"04",X"30",X"02",X"20",X"AD",X"CE",X"00",X"30",X"1E",X"10",X"5F",X"1E",X"10",X"8C",
		X"00",X"00",X"27",X"12",X"30",X"89",X"FF",X"00",X"33",X"C8",X"10",X"11",X"83",X"00",X"30",X"23",
		X"EE",X"CE",X"00",X"10",X"20",X"E9",X"33",X"41",X"47",X"25",X"05",X"57",X"25",X"02",X"20",X"F6",
		X"1F",X"30",X"86",X"01",X"B7",X"C9",X"00",X"10",X"CE",X"F1",X"8D",X"20",X"52",X"86",X"BF",X"1F",
		X"8B",X"1F",X"A8",X"43",X"10",X"CE",X"BF",X"00",X"BD",X"37",X"BC",X"85",X"C0",X"26",X"0A",X"86",
		X"05",X"8E",X"30",X"70",X"C6",X"22",X"BD",X"46",X"23",X"86",X"07",X"8E",X"40",X"90",X"C6",X"22",
		X"BD",X"46",X"23",X"1F",X"30",X"1F",X"98",X"C6",X"22",X"BD",X"46",X"26",X"1F",X"A8",X"85",X"40",
		X"26",X"03",X"7E",X"F8",X"EE",X"10",X"8E",X"FF",X"97",X"86",X"20",X"8E",X"58",X"00",X"30",X"1F",
		X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"00",X"00",X"26",X"F4",X"4A",X"26",X"EE",X"6E",X"A4",X"1F",
		X"03",X"86",X"02",X"1F",X"8B",X"1F",X"30",X"10",X"8E",X"F1",X"EE",X"7E",X"F2",X"69",X"86",X"02",
		X"10",X"8E",X"F1",X"F6",X"20",X"D5",X"10",X"8E",X"F1",X"FC",X"20",X"5D",X"86",X"01",X"10",X"8E",
		X"F2",X"04",X"20",X"C7",X"1F",X"30",X"1F",X"98",X"44",X"44",X"44",X"44",X"10",X"8E",X"F2",X"12",
		X"20",X"57",X"86",X"02",X"10",X"8E",X"F2",X"1A",X"20",X"B1",X"10",X"8E",X"F2",X"20",X"20",X"39",
		X"86",X"01",X"10",X"8E",X"F2",X"28",X"20",X"A3",X"1F",X"30",X"1F",X"98",X"10",X"8E",X"F2",X"32",
		X"20",X"37",X"86",X"02",X"10",X"8E",X"F2",X"3A",X"20",X"91",X"10",X"8E",X"F2",X"40",X"20",X"19",
		X"86",X"05",X"10",X"8E",X"F2",X"48",X"20",X"83",X"1F",X"B8",X"4A",X"1F",X"8B",X"26",X"96",X"10",
		X"8E",X"F2",X"55",X"20",X"04",X"1F",X"30",X"6E",X"E4",X"86",X"3C",X"B7",X"C8",X"0D",X"4C",X"B7",
		X"C8",X"0F",X"86",X"C0",X"B7",X"C8",X"0E",X"6E",X"A4",X"1F",X"89",X"46",X"46",X"46",X"84",X"C0",
		X"B7",X"C8",X"0E",X"86",X"34",X"C5",X"04",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0F",X"86",X"34",
		X"C5",X"08",X"27",X"02",X"86",X"3C",X"B7",X"C8",X"0D",X"6E",X"A4",X"1A",X"3F",X"8E",X"F3",X"1D",
		X"8C",X"F3",X"3D",X"26",X"02",X"6E",X"A4",X"A6",X"01",X"27",X"18",X"A6",X"84",X"5F",X"1F",X"03",
		X"86",X"39",X"EB",X"C0",X"B7",X"CB",X"FF",X"1E",X"03",X"A1",X"02",X"1E",X"03",X"26",X"F3",X"E1",
		X"01",X"26",X"04",X"30",X"02",X"20",X"D9",X"A6",X"84",X"44",X"44",X"44",X"44",X"81",X"0D",X"25",
		X"02",X"80",X"04",X"8B",X"01",X"19",X"1F",X"89",X"86",X"02",X"10",X"CE",X"F2",X"D1",X"7E",X"F1",
		X"DF",X"86",X"BF",X"1F",X"8B",X"86",X"39",X"B7",X"CB",X"FF",X"10",X"CE",X"BF",X"00",X"BD",X"37",
		X"BC",X"1F",X"A8",X"43",X"F7",X"BF",X"15",X"85",X"C0",X"26",X"0A",X"86",X"05",X"8E",X"30",X"70",
		X"C6",X"22",X"BD",X"46",X"23",X"86",X"08",X"8E",X"40",X"90",X"C6",X"22",X"BD",X"46",X"23",X"B6",
		X"BF",X"15",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"C6",X"22",X"BD",X"46",X"26",X"1F",X"A9",X"C5",
		X"40",X"26",X"03",X"7E",X"F8",X"F3",X"10",X"8E",X"FF",X"97",X"7E",X"F1",X"C9",X"00",X"20",X"10",
		X"FC",X"20",X"45",X"30",X"66",X"40",X"B6",X"50",X"11",X"60",X"FD",X"70",X"19",X"80",X"DB",X"90",
		X"00",X"A0",X"00",X"B0",X"00",X"C0",X"00",X"D0",X"6C",X"E0",X"14",X"F0",X"77",X"00",X"63",X"86",
		X"04",X"B7",X"C8",X"05",X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"86",X"FF",X"B7",
		X"BF",X"18",X"BD",X"F4",X"5B",X"B6",X"C8",X"0C",X"46",X"10",X"25",X"06",X"0F",X"BD",X"37",X"BC",
		X"1A",X"BF",X"10",X"8E",X"F3",X"69",X"7E",X"F2",X"59",X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",
		X"0C",X"85",X"02",X"26",X"F4",X"10",X"8E",X"F3",X"7C",X"7E",X"F2",X"8B",X"86",X"BF",X"1F",X"8B",
		X"BD",X"37",X"BC",X"86",X"00",X"BD",X"46",X"32",X"C6",X"03",X"8E",X"70",X"00",X"86",X"39",X"B7",
		X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"16",X"30",X"1F",X"8C",X"00",X"00",X"26",X"ED",
		X"5A",X"26",X"E7",X"10",X"8E",X"F3",X"AF",X"8E",X"00",X"00",X"86",X"FF",X"7E",X"F0",X"9F",X"86",
		X"01",X"B7",X"C9",X"00",X"86",X"BF",X"1F",X"8B",X"BD",X"37",X"BC",X"86",X"01",X"BD",X"46",X"32",
		X"86",X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F4",X"8E",X"9C",X"00",X"6F",
		X"80",X"C6",X"39",X"F7",X"CB",X"FF",X"8C",X"BF",X"01",X"26",X"F4",X"CC",X"A5",X"5A",X"FD",X"BF",
		X"1A",X"B7",X"BF",X"18",X"8D",X"68",X"BD",X"F9",X"2C",X"BD",X"FE",X"BC",X"86",X"02",X"24",X"24",
		X"C6",X"2F",X"8C",X"CD",X"00",X"22",X"02",X"C6",X"1F",X"10",X"CE",X"F4",X"02",X"86",X"03",X"7E",
		X"F1",X"DF",X"10",X"CE",X"BF",X"00",X"8D",X"46",X"86",X"BF",X"1F",X"8B",X"86",X"03",X"C1",X"1F",
		X"22",X"02",X"86",X"04",X"BD",X"37",X"BC",X"BD",X"46",X"32",X"BD",X"F9",X"2C",X"7F",X"BF",X"17",
		X"BD",X"FE",X"3C",X"BD",X"FE",X"46",X"BD",X"F9",X"4F",X"24",X"F8",X"86",X"3F",X"B7",X"C8",X"0E",
		X"4F",X"BD",X"F9",X"5C",X"4F",X"B7",X"C8",X"0E",X"BD",X"F9",X"2C",X"BD",X"F7",X"7D",X"BD",X"F9",
		X"2C",X"BD",X"F6",X"E1",X"BD",X"F9",X"4F",X"24",X"03",X"BD",X"F9",X"2C",X"20",X"75",X"7F",X"C8",
		X"0E",X"86",X"34",X"B7",X"C8",X"0D",X"4C",X"B7",X"C8",X"0F",X"39",X"8E",X"F0",X"12",X"10",X"8E",
		X"C0",X"00",X"EC",X"81",X"ED",X"A1",X"8C",X"F0",X"22",X"25",X"F7",X"39",X"86",X"3C",X"B7",X"C8",
		X"05",X"B7",X"C8",X"07",X"B7",X"C8",X"0D",X"B7",X"C8",X"0F",X"86",X"3F",X"1F",X"8A",X"86",X"8F",
		X"BE",X"C5",X"10",X"30",X"89",X"12",X"34",X"10",X"8E",X"F4",X"8E",X"7E",X"F0",X"9F",X"10",X"8E",
		X"F4",X"95",X"7E",X"F2",X"8B",X"86",X"BF",X"1F",X"8B",X"10",X"CE",X"BF",X"00",X"BD",X"FE",X"BC",
		X"24",X"16",X"86",X"04",X"8C",X"CD",X"00",X"23",X"02",X"86",X"03",X"BD",X"37",X"BC",X"BD",X"46",
		X"32",X"86",X"39",X"B7",X"CB",X"FF",X"20",X"F9",X"8D",X"31",X"10",X"8E",X"F4",X"6C",X"86",X"04",
		X"7E",X"F1",X"CB",X"8D",X"78",X"BD",X"F9",X"2C",X"BD",X"37",X"BC",X"86",X"07",X"B7",X"C0",X"00",
		X"BD",X"F9",X"2C",X"86",X"38",X"B7",X"C0",X"00",X"BD",X"F9",X"2C",X"86",X"C0",X"B7",X"C0",X"00",
		X"BD",X"F9",X"2C",X"8D",X"06",X"BD",X"F9",X"2C",X"7E",X"F9",X"6C",X"8E",X"C0",X"00",X"10",X"8E",
		X"F5",X"2D",X"EC",X"A1",X"ED",X"81",X"86",X"39",X"B7",X"CB",X"FF",X"8C",X"C0",X"10",X"25",X"F2",
		X"CC",X"00",X"00",X"8E",X"00",X"00",X"BF",X"BF",X"15",X"30",X"89",X"0F",X"00",X"ED",X"83",X"34",
		X"02",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"02",X"BC",X"BF",X"15",X"26",X"F0",X"30",X"89",X"09",
		X"00",X"4D",X"26",X"03",X"8E",X"0D",X"00",X"C3",X"11",X"11",X"24",X"DA",X"39",X"05",X"05",X"28",
		X"28",X"80",X"80",X"00",X"00",X"AD",X"AD",X"2D",X"2D",X"A8",X"A8",X"85",X"85",X"BD",X"37",X"BC",
		X"4F",X"BD",X"F7",X"72",X"7F",X"C9",X"00",X"86",X"FF",X"B7",X"C0",X"01",X"86",X"C0",X"B7",X"C0",
		X"02",X"86",X"38",X"B7",X"C0",X"03",X"86",X"07",X"B7",X"C0",X"04",X"10",X"8E",X"F6",X"69",X"CC",
		X"01",X"01",X"AE",X"A4",X"C6",X"39",X"F7",X"CB",X"FF",X"C6",X"01",X"ED",X"81",X"AC",X"22",X"26",
		X"FA",X"31",X"24",X"10",X"8C",X"F6",X"91",X"26",X"E9",X"86",X"11",X"10",X"8E",X"F6",X"49",X"AE",
		X"A4",X"BF",X"BF",X"15",X"A7",X"84",X"7C",X"BF",X"15",X"C6",X"39",X"F7",X"CB",X"FF",X"BE",X"BF",
		X"15",X"AC",X"22",X"26",X"EF",X"31",X"24",X"10",X"8C",X"F6",X"69",X"26",X"E2",X"10",X"8E",X"F6",
		X"91",X"AE",X"A4",X"BF",X"BF",X"15",X"A6",X"24",X"A7",X"84",X"7C",X"BF",X"15",X"C6",X"39",X"F7",
		X"CB",X"FF",X"BE",X"BF",X"15",X"AC",X"22",X"26",X"EF",X"31",X"25",X"10",X"8C",X"F6",X"CD",X"26",
		X"E0",X"10",X"8E",X"F6",X"CD",X"AE",X"A4",X"A6",X"24",X"A7",X"80",X"C6",X"39",X"F7",X"CB",X"FF",
		X"AC",X"22",X"26",X"F5",X"31",X"25",X"10",X"8C",X"F6",X"E1",X"26",X"E9",X"86",X"21",X"B7",X"43",
		X"7E",X"86",X"20",X"B7",X"93",X"7E",X"8E",X"4B",X"0A",X"A6",X"84",X"84",X"F0",X"8A",X"02",X"C6",
		X"39",X"F7",X"CB",X"FF",X"A7",X"80",X"8C",X"4B",X"6D",X"26",X"EE",X"8E",X"4B",X"90",X"A6",X"84",
		X"84",X"F0",X"8A",X"02",X"C6",X"39",X"F7",X"CB",X"FF",X"A7",X"80",X"8C",X"4B",X"F3",X"26",X"EE",
		X"8E",X"0B",X"18",X"BF",X"BF",X"15",X"BE",X"BF",X"15",X"A6",X"84",X"84",X"F0",X"8A",X"01",X"A7",
		X"84",X"F6",X"BF",X"16",X"CB",X"22",X"25",X"05",X"F7",X"BF",X"16",X"20",X"E9",X"C6",X"18",X"F7",
		X"BF",X"16",X"F6",X"BF",X"15",X"CB",X"10",X"F7",X"BF",X"15",X"C1",X"9B",X"26",X"D8",X"C6",X"01",
		X"F7",X"C9",X"00",X"C6",X"39",X"F7",X"CB",X"FF",X"39",X"04",X"07",X"94",X"07",X"04",X"29",X"94",
		X"29",X"04",X"4B",X"94",X"4B",X"04",X"6D",X"94",X"6D",X"04",X"8F",X"94",X"8F",X"04",X"B1",X"94",
		X"B1",X"04",X"D3",X"94",X"D3",X"04",X"F5",X"94",X"F5",X"03",X"07",X"03",X"F5",X"13",X"07",X"13",
		X"F5",X"23",X"07",X"23",X"F5",X"33",X"07",X"33",X"F5",X"43",X"07",X"43",X"F5",X"53",X"07",X"53",
		X"F5",X"63",X"07",X"63",X"F5",X"73",X"07",X"73",X"F5",X"83",X"07",X"83",X"F5",X"93",X"07",X"93",
		X"F5",X"45",X"05",X"52",X"05",X"44",X"45",X"06",X"52",X"06",X"44",X"45",X"07",X"52",X"07",X"00",
		X"45",X"08",X"52",X"08",X"33",X"45",X"09",X"52",X"09",X"33",X"45",X"F3",X"52",X"F3",X"33",X"45",
		X"F4",X"52",X"F4",X"33",X"45",X"F5",X"52",X"F5",X"00",X"45",X"F6",X"52",X"F6",X"44",X"45",X"F7",
		X"52",X"F7",X"44",X"04",X"7E",X"43",X"7E",X"22",X"54",X"7E",X"93",X"7E",X"22",X"02",X"6F",X"02",
		X"8E",X"04",X"03",X"6F",X"03",X"8E",X"30",X"93",X"6F",X"93",X"8E",X"00",X"94",X"6F",X"94",X"8E",
		X"34",X"BD",X"37",X"BC",X"86",X"05",X"BD",X"46",X"32",X"86",X"80",X"B7",X"BF",X"37",X"4F",X"BD",
		X"F9",X"5C",X"BD",X"F9",X"4F",X"25",X"33",X"7A",X"BF",X"37",X"26",X"F2",X"B6",X"F7",X"5A",X"8D",
		X"71",X"8D",X"28",X"8E",X"F7",X"5A",X"A6",X"80",X"BF",X"BF",X"15",X"8D",X"65",X"86",X"80",X"B7",
		X"BF",X"37",X"4F",X"BD",X"F9",X"5C",X"BD",X"F9",X"4F",X"25",X"0F",X"7A",X"BF",X"37",X"26",X"F2",
		X"BE",X"BF",X"15",X"8C",X"F7",X"62",X"25",X"DE",X"20",X"D9",X"39",X"8E",X"00",X"00",X"10",X"8E",
		X"F7",X"62",X"BF",X"BF",X"15",X"30",X"89",X"0F",X"00",X"A6",X"A0",X"1F",X"89",X"ED",X"83",X"C6",
		X"39",X"F7",X"CB",X"FF",X"BC",X"BF",X"15",X"26",X"F2",X"30",X"89",X"09",X"00",X"4D",X"26",X"03",
		X"8E",X"0D",X"00",X"10",X"8C",X"F7",X"72",X"26",X"D9",X"39",X"02",X"03",X"04",X"10",X"18",X"20",
		X"40",X"80",X"00",X"FF",X"11",X"EE",X"22",X"DD",X"33",X"CC",X"44",X"BB",X"55",X"AA",X"66",X"99",
		X"77",X"88",X"8E",X"C0",X"00",X"A7",X"80",X"8C",X"C0",X"10",X"25",X"F9",X"39",X"86",X"0A",X"B7",
		X"BF",X"15",X"BD",X"37",X"BC",X"86",X"06",X"BD",X"46",X"32",X"C6",X"39",X"F7",X"CB",X"FF",X"CE",
		X"BF",X"37",X"6F",X"C0",X"11",X"83",X"BF",X"40",X"23",X"F8",X"CE",X"F8",X"5E",X"8D",X"29",X"86",
		X"34",X"B7",X"C8",X"07",X"C6",X"39",X"F7",X"CB",X"FF",X"8D",X"1D",X"86",X"3C",X"B7",X"C8",X"07",
		X"8D",X"26",X"BD",X"F9",X"4F",X"24",X"0A",X"C6",X"39",X"F7",X"CB",X"FF",X"7A",X"BF",X"15",X"27",
		X"06",X"4F",X"BD",X"F9",X"5C",X"20",X"D3",X"39",X"AE",X"C1",X"27",X"0B",X"10",X"AE",X"C1",X"A6",
		X"84",X"A8",X"A4",X"A7",X"21",X"20",X"F1",X"39",X"CE",X"F8",X"76",X"10",X"8E",X"BF",X"37",X"C6",
		X"01",X"E5",X"21",X"27",X"02",X"8D",X"15",X"33",X"43",X"58",X"24",X"F5",X"C6",X"39",X"F7",X"CB",
		X"FF",X"31",X"22",X"10",X"8C",X"BF",X"40",X"22",X"02",X"20",X"E4",X"39",X"34",X"14",X"86",X"3F",
		X"B7",X"C8",X"0E",X"E8",X"A4",X"E7",X"A4",X"E6",X"E4",X"E5",X"A4",X"26",X"2A",X"E6",X"42",X"27",
		X"4B",X"86",X"40",X"1F",X"01",X"C6",X"39",X"F7",X"CB",X"FF",X"CC",X"40",X"06",X"FD",X"CA",X"06",
		X"BF",X"CA",X"04",X"BF",X"CA",X"04",X"C6",X"00",X"F7",X"CA",X"01",X"C6",X"12",X"F7",X"CA",X"00",
		X"C6",X"39",X"F7",X"CB",X"FF",X"35",X"94",X"E6",X"42",X"27",X"21",X"86",X"40",X"1F",X"01",X"C6",
		X"39",X"F7",X"CB",X"FF",X"C6",X"BB",X"A6",X"C4",X"BD",X"46",X"2C",X"A6",X"41",X"C6",X"39",X"F7",
		X"CB",X"FF",X"C6",X"BB",X"BD",X"46",X"2F",X"86",X"3C",X"B7",X"C8",X"0E",X"35",X"94",X"C8",X"0C",
		X"BF",X"37",X"C8",X"04",X"BF",X"39",X"C8",X"06",X"BF",X"3B",X"00",X"00",X"C8",X"04",X"BF",X"3D",
		X"C8",X"06",X"BF",X"3F",X"00",X"00",X"16",X"FF",X"2C",X"17",X"FF",X"33",X"18",X"FF",X"3A",X"19",
		X"FF",X"41",X"1A",X"FF",X"48",X"1B",X"FF",X"4F",X"1C",X"FF",X"56",X"00",X"00",X"00",X"21",X"F1",
		X"5D",X"6F",X"F1",X"64",X"1F",X"F1",X"6B",X"20",X"F1",X"72",X"1D",X"FF",X"79",X"1E",X"FF",X"80",
		X"72",X"F1",X"87",X"73",X"F1",X"8E",X"70",X"F1",X"95",X"71",X"F1",X"9C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"F2",
		X"A3",X"6F",X"F2",X"AA",X"1F",X"F2",X"B1",X"20",X"F2",X"B8",X"00",X"00",X"00",X"00",X"00",X"00",
		X"72",X"F2",X"BF",X"73",X"F2",X"C6",X"70",X"F2",X"CD",X"71",X"F2",X"D4",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CE",X"F3",
		X"CC",X"20",X"03",X"CE",X"F3",X"A3",X"10",X"CE",X"BF",X"00",X"10",X"8E",X"F9",X"03",X"86",X"01",
		X"7E",X"F1",X"CB",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"10",X"8E",X"F9",X"13",X"86",X"01",
		X"7E",X"F1",X"CB",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F0",X"10",X"8E",X"F9",X"23",X"86",X"01",
		X"7E",X"F1",X"CB",X"B6",X"C8",X"0C",X"85",X"02",X"26",X"F0",X"6E",X"C4",X"B6",X"C8",X"0C",X"85",
		X"02",X"26",X"06",X"86",X"01",X"8D",X"25",X"20",X"F3",X"7F",X"C0",X"00",X"BD",X"37",X"BC",X"20",
		X"07",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"06",X"86",X"01",X"8D",X"10",X"20",X"F3",X"39",X"B6",
		X"C8",X"0C",X"85",X"02",X"27",X"03",X"1A",X"01",X"39",X"1C",X"FE",X"39",X"C6",X"39",X"8E",X"03",
		X"00",X"F7",X"CB",X"FF",X"30",X"1F",X"26",X"F9",X"4A",X"2A",X"F1",X"39",X"86",X"BF",X"1F",X"8B",
		X"BD",X"F4",X"5B",X"8D",X"DA",X"24",X"02",X"8D",X"B3",X"86",X"07",X"BD",X"46",X"32",X"CE",X"CD",
		X"02",X"8E",X"1A",X"30",X"86",X"24",X"34",X"12",X"C6",X"88",X"BD",X"46",X"23",X"1E",X"31",X"BD",
		X"37",X"C2",X"C5",X"F0",X"26",X"08",X"CA",X"F0",X"C5",X"0F",X"26",X"02",X"CA",X"0F",X"1F",X"98",
		X"43",X"34",X"06",X"BD",X"37",X"C5",X"6D",X"E0",X"26",X"12",X"85",X"F0",X"26",X"0E",X"8A",X"F0",
		X"85",X"0F",X"26",X"08",X"8A",X"0F",X"C5",X"F0",X"26",X"02",X"CA",X"F0",X"1F",X"02",X"1E",X"31",
		X"1F",X"10",X"86",X"6A",X"1F",X"01",X"35",X"02",X"C6",X"88",X"BD",X"46",X"26",X"C6",X"39",X"F7",
		X"CB",X"FF",X"1F",X"20",X"34",X"04",X"C6",X"88",X"BD",X"46",X"26",X"35",X"02",X"BD",X"46",X"26",
		X"86",X"39",X"B7",X"CB",X"FF",X"35",X"12",X"30",X"88",X"10",X"4C",X"11",X"83",X"CD",X"38",X"23",
		X"95",X"86",X"2E",X"C6",X"88",X"BD",X"46",X"23",X"1F",X"10",X"86",X"6E",X"1F",X"01",X"1E",X"31",
		X"8E",X"CD",X"20",X"BD",X"37",X"C2",X"F7",X"BF",X"1F",X"BD",X"37",X"C5",X"FD",X"BF",X"20",X"8E",
		X"CD",X"38",X"BD",X"37",X"C2",X"F7",X"BF",X"22",X"BD",X"37",X"C5",X"FD",X"BF",X"23",X"1E",X"31",
		X"8D",X"2C",X"C6",X"88",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"BD",X"46",X"26",X"34",X"10",X"30",
		X"1C",X"86",X"2D",X"BD",X"46",X"20",X"35",X"10",X"86",X"2D",X"BD",X"46",X"20",X"B6",X"BF",X"21",
		X"BD",X"46",X"26",X"86",X"39",X"B7",X"CB",X"FF",X"BD",X"F9",X"2C",X"7E",X"FB",X"4F",X"34",X"30",
		X"8D",X"7A",X"FC",X"BF",X"1F",X"27",X"0F",X"86",X"99",X"34",X"02",X"B7",X"BF",X"21",X"7F",X"BF",
		X"20",X"7F",X"BF",X"1F",X"20",X"4C",X"B6",X"BF",X"21",X"34",X"02",X"FC",X"BF",X"1C",X"FD",X"BF",
		X"1F",X"B6",X"BF",X"1E",X"B7",X"BF",X"21",X"CC",X"00",X"00",X"FD",X"BF",X"1C",X"B7",X"BF",X"1E",
		X"86",X"04",X"78",X"BF",X"21",X"79",X"BF",X"20",X"79",X"BF",X"1F",X"79",X"BF",X"1E",X"4A",X"26",
		X"F1",X"8E",X"BF",X"22",X"10",X"8E",X"BF",X"22",X"CE",X"BF",X"22",X"8D",X"17",X"FC",X"BF",X"1E",
		X"FD",X"BF",X"25",X"FC",X"BF",X"20",X"FD",X"BF",X"27",X"8E",X"BF",X"29",X"8D",X"06",X"8D",X"04",
		X"8D",X"23",X"35",X"B2",X"34",X"70",X"C6",X"04",X"20",X"04",X"34",X"70",X"C6",X"03",X"1C",X"FE",
		X"A6",X"82",X"A9",X"A2",X"19",X"A7",X"C2",X"5A",X"26",X"F6",X"35",X"F0",X"CC",X"00",X"00",X"FD",
		X"BF",X"1C",X"B7",X"BF",X"1E",X"FC",X"BF",X"22",X"26",X"0F",X"B6",X"BF",X"24",X"26",X"0A",X"CC",
		X"00",X"00",X"FD",X"BF",X"1F",X"B7",X"BF",X"21",X"39",X"86",X"07",X"B7",X"BF",X"25",X"8E",X"BF",
		X"1F",X"10",X"8E",X"BF",X"25",X"CE",X"BF",X"29",X"8D",X"35",X"7A",X"BF",X"25",X"26",X"02",X"20",
		X"2E",X"86",X"04",X"78",X"BF",X"21",X"79",X"BF",X"20",X"79",X"BF",X"1F",X"79",X"BF",X"1E",X"79",
		X"BF",X"1D",X"79",X"BF",X"1C",X"4A",X"26",X"EB",X"8D",X"A0",X"25",X"02",X"20",X"DC",X"FC",X"BF",
		X"26",X"FD",X"BF",X"1C",X"B6",X"BF",X"28",X"B7",X"BF",X"1E",X"7C",X"BF",X"21",X"20",X"E9",X"34",
		X"20",X"C6",X"03",X"86",X"99",X"A0",X"A2",X"A7",X"A4",X"5A",X"26",X"F7",X"10",X"AE",X"E4",X"C6",
		X"03",X"1A",X"01",X"A6",X"3F",X"89",X"00",X"19",X"A7",X"A2",X"5A",X"26",X"F6",X"35",X"A0",X"8E",
		X"CC",X"18",X"6F",X"80",X"8C",X"CC",X"23",X"25",X"F9",X"BD",X"37",X"BC",X"BD",X"F9",X"4F",X"24",
		X"03",X"BD",X"F9",X"2C",X"86",X"08",X"BD",X"46",X"32",X"CE",X"CC",X"00",X"8E",X"1A",X"20",X"86",
		X"30",X"34",X"12",X"C6",X"22",X"BD",X"46",X"2C",X"F7",X"BF",X"29",X"F7",X"BF",X"1C",X"1F",X"12",
		X"BD",X"FD",X"2A",X"33",X"42",X"C6",X"39",X"F7",X"CB",X"FF",X"35",X"12",X"30",X"0A",X"4C",X"11",
		X"83",X"CC",X"24",X"2D",X"DC",X"86",X"09",X"BD",X"46",X"35",X"7F",X"BF",X"1C",X"4F",X"F6",X"BF",
		X"29",X"8E",X"6E",X"34",X"BD",X"46",X"2C",X"B6",X"CC",X"07",X"84",X"0F",X"81",X"09",X"26",X"08",
		X"86",X"5D",X"8E",X"70",X"3E",X"BD",X"46",X"2C",X"10",X"8E",X"16",X"20",X"CE",X"CC",X"00",X"1F",
		X"21",X"86",X"2E",X"C6",X"33",X"FD",X"BF",X"37",X"BD",X"46",X"29",X"86",X"39",X"B7",X"CB",X"FF",
		X"B6",X"C8",X"04",X"84",X"03",X"27",X"02",X"8D",X"1A",X"B6",X"C8",X"04",X"84",X"C0",X"27",X"03",
		X"BD",X"FC",X"86",X"C6",X"3C",X"F7",X"C8",X"07",X"BD",X"F9",X"4F",X"24",X"DE",X"BD",X"F9",X"2C",
		X"7E",X"37",X"B0",X"B7",X"BF",X"3B",X"B1",X"BF",X"39",X"27",X"15",X"7F",X"BF",X"3A",X"B6",X"BF",
		X"3B",X"B7",X"BF",X"39",X"86",X"02",X"BD",X"F9",X"5C",X"B6",X"C8",X"04",X"84",X"03",X"26",X"1D",
		X"C6",X"05",X"F7",X"BF",X"3C",X"B6",X"C8",X"04",X"84",X"03",X"26",X"04",X"7F",X"BF",X"39",X"39",
		X"86",X"02",X"BD",X"F9",X"5C",X"7A",X"BF",X"3C",X"26",X"EB",X"B6",X"C8",X"04",X"85",X"02",X"26",
		X"22",X"85",X"01",X"27",X"42",X"10",X"8C",X"16",X"20",X"27",X"3C",X"8D",X"3F",X"31",X"36",X"33",
		X"5E",X"11",X"83",X"CC",X"12",X"26",X"0A",X"7D",X"BF",X"19",X"27",X"05",X"31",X"A8",X"C4",X"33",
		X"54",X"20",X"1C",X"10",X"8C",X"16",X"CA",X"27",X"1E",X"8D",X"21",X"31",X"2A",X"33",X"42",X"11",
		X"83",X"CC",X"08",X"26",X"0A",X"7D",X"BF",X"19",X"27",X"05",X"31",X"A8",X"3C",X"33",X"4C",X"1F",
		X"21",X"FC",X"BF",X"37",X"BD",X"46",X"29",X"4F",X"BD",X"F9",X"5C",X"39",X"1F",X"21",X"B6",X"BF",
		X"37",X"5F",X"BD",X"46",X"29",X"39",X"B7",X"BF",X"3B",X"B1",X"BF",X"3D",X"27",X"15",X"7F",X"BF",
		X"3E",X"B6",X"BF",X"3B",X"B7",X"BF",X"3D",X"86",X"02",X"BD",X"F9",X"5C",X"B6",X"C8",X"04",X"84",
		X"C0",X"26",X"1E",X"C6",X"08",X"F7",X"BF",X"40",X"B6",X"C8",X"04",X"84",X"C0",X"26",X"04",X"7F",
		X"BF",X"3E",X"39",X"4F",X"BD",X"F9",X"5C",X"7A",X"BF",X"40",X"26",X"EC",X"B6",X"C8",X"04",X"84",
		X"C0",X"34",X"02",X"1F",X"31",X"BD",X"37",X"BF",X"34",X"02",X"5F",X"F7",X"BF",X"29",X"8D",X"5A",
		X"C6",X"39",X"F7",X"CB",X"FF",X"8E",X"FD",X"06",X"1F",X"30",X"30",X"85",X"35",X"06",X"C5",X"40",
		X"26",X"0C",X"C5",X"80",X"27",X"14",X"A1",X"84",X"27",X"10",X"8B",X"99",X"20",X"06",X"A1",X"01",
		X"27",X"08",X"8B",X"01",X"19",X"1F",X"31",X"BD",X"37",X"C8",X"C6",X"22",X"F7",X"BF",X"29",X"BD",
		X"FD",X"2A",X"4F",X"7E",X"F9",X"5C",X"15",X"99",X"01",X"79",X"00",X"99",X"00",X"09",X"00",X"99",
		X"00",X"99",X"00",X"99",X"01",X"99",X"00",X"99",X"00",X"99",X"00",X"09",X"03",X"20",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"1F",X"30",X"54",X"8E",X"FD",X"7E",
		X"30",X"85",X"6D",X"84",X"2B",X"2C",X"1F",X"31",X"BD",X"37",X"BF",X"11",X"83",X"CC",X"06",X"26",
		X"0A",X"B7",X"BF",X"19",X"7D",X"BF",X"1C",X"26",X"02",X"8D",X"45",X"85",X"F0",X"26",X"02",X"8A",
		X"F0",X"34",X"02",X"1F",X"20",X"86",X"6A",X"1F",X"01",X"35",X"02",X"F6",X"BF",X"29",X"BD",X"46",
		X"2F",X"39",X"1F",X"31",X"BD",X"37",X"C2",X"86",X"0D",X"5D",X"27",X"02",X"86",X"44",X"34",X"02",
		X"1F",X"20",X"86",X"6A",X"1F",X"01",X"35",X"02",X"F6",X"BF",X"29",X"7E",X"46",X"2C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",
		X"34",X"76",X"8E",X"04",X"38",X"BF",X"CA",X"06",X"8E",X"6A",X"48",X"BF",X"CA",X"04",X"5F",X"F7",
		X"CA",X"01",X"C6",X"12",X"F7",X"CA",X"00",X"8E",X"FE",X"00",X"81",X"09",X"26",X"0F",X"34",X"12",
		X"86",X"5D",X"F6",X"BF",X"29",X"8E",X"70",X"3E",X"BD",X"46",X"2C",X"35",X"12",X"1F",X"89",X"58",
		X"34",X"04",X"58",X"EB",X"E0",X"3A",X"33",X"42",X"1E",X"31",X"8C",X"CC",X"14",X"27",X"2F",X"A6",
		X"C0",X"BD",X"37",X"C8",X"C6",X"39",X"F7",X"CB",X"FF",X"1E",X"31",X"31",X"2A",X"34",X"10",X"30",
		X"5E",X"BD",X"37",X"BF",X"85",X"F0",X"26",X"02",X"8A",X"F0",X"34",X"02",X"1F",X"20",X"86",X"6A",
		X"1F",X"01",X"35",X"02",X"F6",X"BF",X"29",X"BD",X"46",X"2F",X"35",X"10",X"20",X"CA",X"35",X"F6",
		X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"04",X"01",X"02",X"04",X"00",X"06",X"00",X"01",X"01",
		X"00",X"00",X"01",X"04",X"01",X"01",X"00",X"00",X"01",X"16",X"06",X"02",X"00",X"00",X"01",X"04",
		X"01",X"02",X"00",X"00",X"01",X"00",X"04",X"01",X"00",X"00",X"01",X"00",X"02",X"01",X"00",X"00",
		X"01",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"37",X"BC",X"CC",
		X"FE",X"01",X"FD",X"BF",X"38",X"39",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",X"F9",X"5C",
		X"4F",X"B7",X"C8",X"0E",X"86",X"03",X"BD",X"F9",X"5C",X"86",X"3F",X"B7",X"C8",X"0E",X"86",X"03",
		X"BD",X"F9",X"5C",X"FC",X"BF",X"38",X"84",X"3F",X"B7",X"C8",X"0E",X"C6",X"99",X"8E",X"3A",X"80",
		X"86",X"22",X"BD",X"46",X"23",X"B6",X"BF",X"39",X"8A",X"F0",X"C6",X"99",X"BD",X"46",X"26",X"86",
		X"40",X"B7",X"BF",X"37",X"86",X"01",X"BD",X"F9",X"5C",X"BD",X"F9",X"4F",X"25",X"05",X"7A",X"BF",
		X"37",X"26",X"F1",X"B6",X"BF",X"17",X"26",X"06",X"B6",X"C8",X"0C",X"46",X"24",X"1D",X"8E",X"57",
		X"80",X"B6",X"BF",X"39",X"8A",X"F0",X"C6",X"00",X"BD",X"46",X"26",X"FC",X"BF",X"38",X"1A",X"01",
		X"49",X"5C",X"C1",X"07",X"25",X"02",X"8D",X"87",X"FD",X"BF",X"38",X"39",X"8E",X"CC",X"00",X"10",
		X"8E",X"9C",X"00",X"A6",X"80",X"A7",X"A0",X"8C",X"D0",X"00",X"26",X"F7",X"C6",X"06",X"FE",X"BF",
		X"1A",X"10",X"BE",X"BF",X"19",X"8E",X"CC",X"00",X"BD",X"FF",X"23",X"A7",X"80",X"86",X"39",X"B7",
		X"CB",X"FF",X"8C",X"D0",X"00",X"26",X"F1",X"10",X"BF",X"BF",X"19",X"FF",X"BF",X"1A",X"8E",X"CC",
		X"00",X"BD",X"FF",X"23",X"A8",X"80",X"84",X"0F",X"26",X"24",X"86",X"39",X"B7",X"CB",X"FF",X"8C",
		X"D0",X"00",X"26",X"ED",X"5A",X"26",X"C7",X"8D",X"03",X"1C",X"FE",X"39",X"CE",X"9C",X"00",X"10",
		X"8E",X"CC",X"00",X"A6",X"C0",X"A7",X"A0",X"10",X"8C",X"D0",X"00",X"26",X"F6",X"39",X"8D",X"EC",
		X"1A",X"01",X"39",X"34",X"04",X"F6",X"BF",X"19",X"86",X"03",X"3D",X"CB",X"11",X"B6",X"BF",X"1B",
		X"44",X"44",X"44",X"B8",X"BF",X"1B",X"44",X"76",X"BF",X"1A",X"76",X"BF",X"1B",X"FB",X"BF",X"1B",
		X"F9",X"BF",X"1A",X"F7",X"BF",X"19",X"B6",X"BF",X"19",X"35",X"84",X"20",X"53",X"50",X"4C",X"41",
		X"54",X"20",X"2D",X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"20",X"28",
		X"43",X"29",X"20",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",X"4C",X"49",X"41",X"4D",X"53",
		X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",X"53",X"20",X"49",X"4E",X"43",
		X"2E",X"20",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",X"20",X"52",X"45",
		X"53",X"45",X"52",X"56",X"45",X"44",X"20",X"BD",X"37",X"F8",X"BD",X"37",X"EC",X"27",X"40",X"86",
		X"39",X"B7",X"CB",X"FF",X"BD",X"37",X"FB",X"86",X"39",X"B7",X"CB",X"FF",X"BD",X"37",X"F5",X"86",
		X"39",X"B7",X"CB",X"FF",X"BD",X"37",X"BC",X"86",X"39",X"B7",X"CB",X"FF",X"BD",X"37",X"F2",X"BD",
		X"37",X"EF",X"BD",X"37",X"E9",X"BD",X"37",X"EC",X"27",X"1A",X"86",X"0B",X"BD",X"46",X"32",X"86",
		X"39",X"B7",X"CB",X"FF",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"F4",X"6E",X"9F",X"EF",X"FE",X"BD",
		X"37",X"E9",X"20",X"F7",X"86",X"0C",X"20",X"E4",X"6E",X"9F",X"EF",X"F8",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"FF",X"E8",X"F0",X"00",X"F0",X"00",X"F0",X"00",
		X"0A",X"6A",X"0A",X"92",X"15",X"C6",X"15",X"EE",X"0C",X"38",X"0E",X"AE",X"11",X"24",X"11",X"4C",
		X"13",X"BC",X"13",X"E4",X"2C",X"D3",X"2C",X"AB",X"17",X"98",X"17",X"70",X"00",X"2B",X"00",X"00",
		X"00",X"00",X"93",X"01",X"00",X"FB",X"01",X"05",X"FE",X"00",X"FD",X"08",X"0A",X"0D",X"1D",X"D3",
		X"00",X"03",X"DD",X"1D",X"00",X"00",X"11",X"DD",X"77",X"7B",X"D1",X"10",X"00",X"00",X"D1",X"1D",
		X"33",X"3D",X"11",X"D0",X"00",X"00",X"D1",X"11",X"D3",X"D1",X"11",X"D0",X"00",X"0D",X"11",X"11",
		X"11",X"11",X"31",X"1D",X"00",X"01",X"C1",X"11",X"11",X"11",X"CD",X"D1",X"00",X"0E",X"7C",X"D1",
		X"11",X"1D",X"74",X"7D",X"00",X"00",X"C4",X"C7",X"74",X"4C",X"C4",X"C0",X"00",X"39",X"7A",X"4C",
		X"00",X"0E",X"4C",X"79",X"30",X"E7",X"77",X"E4",X"C0",X"C4",X"E7",X"77",X"E0",X"01",X"0D",X"02",
		X"0C",X"02",X"0C",X"02",X"0C",X"01",X"0D",X"01",X"0D",X"01",X"0D",X"02",X"0C",X"00",X"0E",X"00",
		X"0E",X"FF",X"FF",X"09",X"0A",X"00",X"D1",X"DD",X"30",X"00",X"3D",X"D1",X"D0",X"00",X"00",X"01",
		X"1D",X"D7",X"77",X"BD",X"11",X"00",X"00",X"00",X"0D",X"11",X"D3",X"33",X"D1",X"1D",X"00",X"00",
		X"00",X"0D",X"11",X"1D",X"3D",X"11",X"1D",X"00",X"00",X"00",X"B1",X"11",X"11",X"11",X"11",X"11",
		X"D0",X"00",X"00",X"DD",X"D3",X"33",X"73",X"33",X"9C",X"D0",X"00",X"00",X"07",X"C9",X"33",X"33",
		X"99",X"C4",X"00",X"00",X"73",X"04",X"4C",X"CC",X"44",X"CC",X"44",X"03",X"70",X"E7",X"E3",X"4C",
		X"00",X"00",X"0C",X"43",X"77",X"E0",X"00",X"E7",X"C4",X"00",X"00",X"04",X"7C",X"E0",X"00",X"02",
		X"0E",X"03",X"0D",X"03",X"0D",X"03",X"0D",X"02",X"0E",X"02",X"0E",X"03",X"0D",X"00",X"10",X"00",
		X"10",X"02",X"0E",X"FF",X"FF",X"0E",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"93",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",
		X"00",X"E3",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"30",X"00",X"3E",X"00",X"00",X"00",X"E7",
		X"E0",X"00",X"00",X"00",X"00",X"00",X"03",X"30",X"0E",X"7E",X"00",X"00",X"00",X"0E",X"7C",X"00",
		X"00",X"00",X"00",X"00",X"03",X"90",X"C7",X"E0",X"00",X"00",X"00",X"0E",X"C4",X"E0",X"00",X"00",
		X"00",X"00",X"B3",X"7E",X"4E",X"E0",X"00",X"03",X"00",X"00",X"C4",X"4E",X"B1",X"DE",X"0E",X"D1",
		X"DD",X"44",X"7C",X"00",X"00",X"73",X"03",X"00",X"0E",X"44",X"CB",X"D1",X"31",X"1D",X"B4",X"CC",
		X"E0",X"00",X"00",X"07",X"33",X"33",X"37",X"C4",X"4C",X"CD",X"DD",X"CC",X"44",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"E7",X"39",X"7C",X"44",X"44",X"44",X"44",X"4C",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EC",X"44",X"C4",X"4C",X"E0",X"00",X"00",X"00",X"00",X"15",X"17",X"15",
		X"16",X"13",X"15",X"14",X"15",X"04",X"19",X"04",X"19",X"05",X"18",X"05",X"18",X"01",X"17",X"00",
		X"16",X"01",X"14",X"04",X"13",X"0A",X"12",X"FF",X"FF",X"01",X"E3",X"00",X"00",X"00",X"02",X"A4",
		X"00",X"00",X"00",X"07",X"15",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"70",
		X"7E",X"00",X"00",X"00",X"00",X"05",X"70",X"00",X"E0",X"00",X"00",X"00",X"E2",X"2E",X"00",X"00",
		X"00",X"00",X"0E",X"21",X"79",X"E0",X"00",X"00",X"00",X"07",X"12",X"92",X"70",X"00",X"00",X"00",
		X"02",X"22",X"27",X"90",X"00",X"00",X"00",X"09",X"12",X"99",X"70",X"00",X"00",X"00",X"09",X"92",
		X"29",X"90",X"00",X"00",X"00",X"09",X"0E",X"70",X"70",X"00",X"00",X"00",X"E2",X"12",X"29",X"2E",
		X"00",X"00",X"5B",X"79",X"02",X"2E",X"97",X"E5",X"00",X"05",X"E9",X"9E",X"09",X"9E",X"50",X"00",
		X"00",X"57",X"92",X"29",X"95",X"00",X"00",X"00",X"57",X"29",X"99",X"75",X"00",X"00",X"00",X"57",
		X"92",X"79",X"75",X"00",X"00",X"00",X"57",X"72",X"99",X"E5",X"00",X"00",X"00",X"05",X"79",X"97",
		X"50",X"00",X"00",X"00",X"00",X"57",X"75",X"00",X"00",X"00",X"00",X"05",X"50",X"05",X"50",X"00",
		X"00",X"07",X"55",X"00",X"00",X"55",X"E0",X"00",X"07",X"07",X"06",X"09",X"05",X"0A",X"04",X"07",
		X"03",X"08",X"03",X"08",X"03",X"08",X"03",X"08",X"03",X"08",X"03",X"08",X"02",X"09",X"00",X"0B",
		X"01",X"0A",X"02",X"09",X"02",X"09",X"02",X"09",X"02",X"09",X"03",X"08",X"04",X"07",X"03",X"08",
		X"01",X"0A",X"FF",X"FF",X"07",X"15",X"00",X"00",X"00",X"09",X"E0",X"E0",X"00",X"00",X"00",X"00",
		X"70",X"0E",X"00",X"00",X"00",X"00",X"05",X"70",X"00",X"00",X"00",X"00",X"00",X"E2",X"2E",X"00",
		X"00",X"00",X"00",X"0E",X"21",X"79",X"E0",X"00",X"00",X"00",X"07",X"12",X"92",X"70",X"00",X"00",
		X"00",X"02",X"22",X"27",X"90",X"00",X"00",X"00",X"09",X"12",X"99",X"70",X"00",X"00",X"00",X"09",
		X"92",X"29",X"90",X"00",X"00",X"00",X"09",X"0E",X"70",X"70",X"00",X"00",X"00",X"E2",X"12",X"29",
		X"2E",X"00",X"00",X"5B",X"79",X"02",X"2E",X"97",X"E5",X"00",X"05",X"E9",X"9E",X"09",X"9E",X"50",
		X"00",X"00",X"57",X"92",X"29",X"95",X"00",X"00",X"00",X"57",X"29",X"99",X"75",X"00",X"00",X"00",
		X"57",X"92",X"79",X"75",X"00",X"00",X"00",X"57",X"72",X"99",X"E5",X"00",X"00",X"00",X"05",X"79",
		X"97",X"50",X"00",X"00",X"00",X"00",X"57",X"75",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",
		X"00",X"00",X"00",X"E5",X"5E",X"05",X"5E",X"00",X"00",X"07",X"0A",X"06",X"09",X"05",X"06",X"04",
		X"07",X"03",X"08",X"03",X"08",X"03",X"08",X"03",X"08",X"03",X"08",X"03",X"08",X"02",X"09",X"00",
		X"0B",X"01",X"0A",X"02",X"09",X"02",X"09",X"02",X"09",X"02",X"09",X"03",X"08",X"04",X"07",X"05",
		X"06",X"02",X"09",X"FF",X"FF",X"03",X"74",X"00",X"00",X"00",X"03",X"D2",X"00",X"80",X"FB",X"04",
		X"44",X"FE",X"00",X"FE",X"07",X"0A",X"AB",X"DE",X"C0",X"00",X"CE",X"DB",X"A0",X"0A",X"AD",X"EC",
		X"CC",X"ED",X"AA",X"00",X"0B",X"BA",X"D4",X"CC",X"DA",X"AB",X"00",X"00",X"BB",X"AD",X"ED",X"AB",
		X"B0",X"00",X"00",X"BB",X"BA",X"DA",X"BB",X"B0",X"00",X"00",X"F6",X"88",X"88",X"88",X"F0",X"00",
		X"00",X"68",X"A0",X"00",X"A8",X"80",X"00",X"00",X"88",X"00",X"00",X"08",X"80",X"00",X"0A",X"D8",
		X"00",X"00",X"08",X"DA",X"00",X"AD",X"DA",X"00",X"00",X"0A",X"DD",X"A0",X"00",X"0C",X"01",X"0B",
		X"01",X"0B",X"02",X"0A",X"02",X"0A",X"02",X"0A",X"02",X"0A",X"02",X"0A",X"01",X"0B",X"00",X"0C",
		X"FF",X"FF",X"08",X"0B",X"0D",X"B0",X"00",X"00",X"00",X"00",X"BD",X"00",X"0A",X"AD",X"CC",X"00",
		X"0C",X"CD",X"AA",X"00",X"00",X"BA",X"DC",X"CC",X"CC",X"DA",X"B0",X"00",X"00",X"BB",X"AB",X"AA",
		X"AB",X"AB",X"B0",X"00",X"00",X"0B",X"BB",X"BA",X"BB",X"BB",X"00",X"00",X"00",X"0F",X"66",X"88",
		X"88",X"8F",X"00",X"00",X"00",X"06",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"F6",X"8F",X"00",
		X"0F",X"86",X"F0",X"00",X"00",X"B8",X"00",X"00",X"00",X"08",X"B0",X"00",X"0A",X"DB",X"00",X"00",
		X"00",X"0B",X"DA",X"00",X"AD",X"B0",X"00",X"00",X"00",X"00",X"DD",X"A0",X"01",X"0D",X"01",X"0D",
		X"02",X"0C",X"02",X"0C",X"03",X"0B",X"03",X"0B",X"03",X"0B",X"02",X"0C",X"02",X"0C",X"01",X"0D",
		X"00",X"0E",X"FF",X"FF",X"0D",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"37",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"70",X"00",X"00",X"00",X"0D",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"AB",X"C0",X"01",X"D0",X"00",X"0A",X"DB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"00",X"BD",X"A0",X"00",X"00",X"AD",X"80",X"00",X"00",X"00",X"00",X"0A",X"BB",X"08",X"DA",
		X"00",X"00",X"00",X"AD",X"A8",X"00",X"B0",X"00",X"00",X"BA",X"BA",X"8A",X"DA",X"00",X"03",X"00",
		X"00",X"66",X"80",X"AD",X"00",X"0D",X"AB",X"B8",X"68",X"00",X"00",X"73",X"07",X"00",X"06",X"88",
		X"AB",X"C7",X"CB",X"BA",X"86",X"80",X"00",X"00",X"07",X"33",X"4B",X"BA",X"68",X"88",X"AA",X"AA",
		X"88",X"68",X"00",X"00",X"00",X"00",X"00",X"CB",X"BB",X"A8",X"88",X"88",X"88",X"88",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F8",X"68",X"86",X"8F",X"00",X"00",X"00",X"00",X"04",
		X"FE",X"00",X"00",X"00",X"05",X"4A",X"FF",X"80",X"F9",X"05",X"96",X"FD",X"80",X"FC",X"06",X"09",
		X"07",X"3C",X"33",X"C3",X"37",X"00",X"03",X"34",X"43",X"9C",X"30",X"00",X"0C",X"C4",X"43",X"34",
		X"40",X"00",X"C4",X"44",X"44",X"44",X"C0",X"00",X"0C",X"44",X"CC",X"E0",X"00",X"00",X"00",X"C4",
		X"4C",X"C0",X"00",X"00",X"00",X"03",X"00",X"30",X"00",X"00",X"00",X"C3",X"00",X"43",X"00",X"C0",
		X"0C",X"4E",X"00",X"40",X"44",X"00",X"01",X"09",X"01",X"08",X"01",X"08",X"00",X"08",X"01",X"06",
		X"02",X"06",X"03",X"06",X"02",X"0A",X"01",X"09",X"FF",X"FF",X"06",X"09",X"00",X"73",X"C3",X"3C",
		X"33",X"70",X"00",X"3C",X"93",X"34",X"73",X"00",X"00",X"44",X"33",X"44",X"CC",X"00",X"00",X"C4",
		X"44",X"44",X"44",X"C0",X"00",X"00",X"EE",X"C4",X"4C",X"00",X"00",X"00",X"CC",X"44",X"C0",X"00",
		X"00",X"00",X"30",X"03",X"00",X"00",X"C0",X"03",X"40",X"03",X"C0",X"00",X"04",X"40",X"C0",X"0E",
		X"4C",X"00",X"02",X"0A",X"02",X"09",X"02",X"09",X"02",X"0A",X"04",X"09",X"04",X"08",X"04",X"07",
		X"00",X"08",X"01",X"09",X"FF",X"FF",X"0D",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"73",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"40",X"00",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"04",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"94",X"00",X"00",X"00",X"E4",X"30",X"00",X"00",X"00",X"00",X"00",X"03",
		X"03",X"4E",X"00",X"00",X"00",X"0C",X"33",X"00",X"00",X"00",X"00",X"00",X"03",X"73",X"C0",X"00",
		X"03",X"00",X"CC",X"73",X"30",X"3C",X"73",X"37",X"C7",X"33",X"37",X"CC",X"00",X"73",X"07",X"00",
		X"0E",X"39",X"CC",X"73",X"97",X"CC",X"33",X"70",X"00",X"00",X"0E",X"93",X"43",X"37",X"73",X"3C",
		X"CC",X"CC",X"C3",X"3E",X"00",X"00",X"00",X"00",X"00",X"CC",X"00",X"0C",X"3C",X"44",X"44",X"C9",
		X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EC",X"44",X"44",X"CE",X"00",X"00",X"00",
		X"00",X"06",X"50",X"00",X"00",X"00",X"06",X"B7",X"01",X"00",X"FC",X"07",X"15",X"FE",X"00",X"FD",
		X"09",X"09",X"00",X"0E",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"72",X"73",X"00",X"00",
		X"03",X"79",X"70",X"00",X"00",X"09",X"97",X"30",X"00",X"37",X"99",X"00",X"00",X"00",X"00",X"72",
		X"27",X"C7",X"29",X"70",X"00",X"00",X"00",X"00",X"E9",X"22",X"22",X"29",X"E0",X"00",X"00",X"00",
		X"00",X"29",X"77",X"97",X"79",X"20",X"00",X"00",X"0D",X"1D",X"D7",X"00",X"00",X"07",X"DD",X"1D",
		X"00",X"B1",X"11",X"6D",X"00",X"00",X"0D",X"61",X"11",X"B0",X"AD",X"DB",X"A0",X"00",X"00",X"00",
		X"AB",X"DD",X"A0",X"03",X"0D",X"02",X"0E",X"03",X"0D",X"04",X"0C",X"04",X"0C",X"04",X"0C",X"01",
		X"0F",X"00",X"10",X"00",X"10",X"FF",X"FF",X"08",X"09",X"07",X"70",X"00",X"00",X"00",X"00",X"77",
		X"00",X"02",X"27",X"30",X"00",X"00",X"37",X"92",X"00",X"00",X"E9",X"73",X"00",X"03",X"79",X"E0",
		X"00",X"00",X"07",X"92",X"7C",X"72",X"97",X"00",X"00",X"00",X"0E",X"92",X"22",X"22",X"9E",X"00",
		X"00",X"00",X"00",X"A9",X"70",X"79",X"A0",X"00",X"00",X"0D",X"1D",X"DA",X"D0",X"DA",X"DD",X"1D",
		X"00",X"B1",X"11",X"DD",X"B0",X"BD",X"D3",X"11",X"B0",X"AD",X"DD",X"BA",X"00",X"0A",X"BD",X"DD",
		X"A0",X"01",X"0D",X"01",X"0D",X"02",X"0C",X"03",X"0B",X"03",X"0B",X"04",X"0A",X"01",X"0D",X"00",
		X"0E",X"00",X"0E",X"FF",X"FF",X"0D",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"70",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"93",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"0D",X"1B",X"00",X"00",X"00",X"00",
		X"00",X"02",X"90",X"B1",X"D0",X"00",X"00",X"01",X"1D",X"00",X"00",X"00",X"00",X"00",X"02",X"90",
		X"D1",X"10",X"00",X"00",X"0B",X"1B",X"70",X"00",X"00",X"00",X"00",X"79",X"79",X"B1",X"B0",X"03",
		X"00",X"00",X"BD",X"27",X"E7",X"70",X"00",X"79",X"97",X"72",X"DB",X"00",X"73",X"03",X"00",X"DD",
		X"92",X"77",X"79",X"C9",X"97",X"79",X"29",X"DD",X"00",X"07",X"33",X"31",X"77",X"79",X"29",X"77",
		X"77",X"79",X"29",X"00",X"00",X"00",X"00",X"00",X"D9",X"99",X"7E",X"79",X"22",X"22",X"22",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"79",X"99",X"97",X"E0",X"00",X"00",X"00",
		X"15",X"17",X"15",X"16",X"13",X"15",X"14",X"15",X"13",X"14",X"05",X"18",X"05",X"18",X"05",X"18",
		X"01",X"17",X"00",X"17",X"01",X"13",X"04",X"12",X"0B",X"12",X"FF",X"FF",X"07",X"E1",X"01",X"00",
		X"FB",X"07",X"07",X"00",X"E4",X"CE",X"E0",X"EC",X"00",X"00",X"0E",X"EC",X"EC",X"73",X"37",X"EC",
		X"00",X"7C",X"E3",X"33",X"33",X"33",X"E9",X"70",X"37",X"37",X"07",X"27",X"07",X"37",X"30",X"0E",
		X"33",X"9E",X"CE",X"93",X"3E",X"00",X"00",X"73",X"EC",X"CE",X"E3",X"70",X"00",X"00",X"00",X"03",
		X"33",X"00",X"00",X"00",X"02",X"09",X"01",X"0B",X"00",X"0C",X"00",X"0C",X"01",X"0B",X"02",X"0A",
		X"05",X"07",X"FF",X"FF",X"08",X"29",X"00",X"80",X"FB",X"07",X"07",X"00",X"EE",X"CE",X"EE",X"0E",
		X"00",X"00",X"0E",X"73",X"39",X"EE",X"33",X"EE",X"00",X"EC",X"93",X"23",X"33",X"23",X"9C",X"E0",
		X"3E",X"37",X"07",X"97",X"07",X"3E",X"30",X"77",X"39",X"93",X"23",X"99",X"37",X"70",X"00",X"73",
		X"3E",X"73",X"33",X"70",X"00",X"00",X"00",X"09",X"37",X"00",X"00",X"00",X"02",X"09",X"01",X"0B",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"02",X"0A",X"05",X"07",X"FF",X"FF",X"08",X"71",X"FF",X"80",
		X"F9",X"07",X"07",X"00",X"07",X"92",X"97",X"E9",X"E0",X"00",X"00",X"72",X"92",X"99",X"33",X"9E",
		X"00",X"00",X"29",X"00",X"39",X"00",X"92",X"00",X"E9",X"27",X"43",X"32",X"34",X"99",X"70",X"22",
		X"77",X"33",X"4C",X"33",X"72",X"20",X"99",X"97",X"93",X"33",X"39",X"E2",X"90",X"09",X"29",X"0E",
		X"37",X"07",X"29",X"00",X"03",X"0A",X"02",X"0B",X"02",X"0B",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"01",X"0B",X"FF",X"FF",X"08",X"B9",X"01",X"00",X"FC",X"07",X"07",X"00",X"EC",X"91",X"73",X"9C",
		X"E0",X"00",X"3C",X"E7",X"39",X"39",X"37",X"EC",X"30",X"3E",X"73",X"70",X"70",X"73",X"7E",X"30",
		X"03",X"34",X"33",X"23",X"34",X"33",X"00",X"00",X"33",X"E0",X"D0",X"E3",X"30",X"00",X"00",X"00",
		X"3E",X"0E",X"30",X"00",X"00",X"00",X"00",X"03",X"33",X"00",X"00",X"00",X"02",X"0A",X"00",X"0C",
		X"00",X"0C",X"01",X"0B",X"02",X"0A",X"04",X"08",X"05",X"07",X"FF",X"FF",X"09",X"01",X"FC",X"00",
		X"01",X"06",X"04",X"00",X"00",X"00",X"00",X"D1",X"10",X"33",X"70",X"03",X"00",X"71",X"10",X"0E",
		X"33",X"33",X"93",X"39",X"D0",X"00",X"00",X"07",X"33",X"37",X"00",X"08",X"0A",X"00",X"0A",X"01",
		X"0A",X"05",X"09",X"FF",X"FF",X"09",X"2A",X"07",X"00",X"01",X"06",X"04",X"11",X"D0",X"00",X"00",
		X"00",X"00",X"11",X"70",X"03",X"00",X"73",X"30",X"D9",X"33",X"93",X"33",X"3E",X"00",X"07",X"33",
		X"37",X"00",X"00",X"00",X"00",X"02",X"00",X"0A",X"00",X"09",X"01",X"05",X"FF",X"FF",X"09",X"53",
		X"FC",X"00",X"00",X"06",X"03",X"33",X"70",X"03",X"00",X"00",X"70",X"0E",X"33",X"33",X"43",X"33",
		X"30",X"00",X"00",X"0C",X"00",X"70",X"00",X"00",X"0A",X"01",X"0A",X"05",X"08",X"FF",X"FF",X"09",
		X"74",X"04",X"80",X"00",X"06",X"03",X"3E",X"00",X"03",X"00",X"73",X"30",X"33",X"33",X"43",X"33",
		X"3E",X"00",X"00",X"70",X"0C",X"00",X"00",X"00",X"00",X"0A",X"00",X"09",X"02",X"05",X"FF",X"FF",
		X"09",X"95",X"FB",X"00",X"01",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"B0",X"33",X"70",X"03",
		X"00",X"0B",X"B0",X"0E",X"33",X"33",X"CD",X"BB",X"B0",X"00",X"00",X"07",X"CA",X"BA",X"00",X"0A",
		X"0A",X"00",X"0A",X"01",X"0A",X"05",X"09",X"FF",X"FF",X"09",X"BE",X"05",X"80",X"01",X"06",X"04",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"03",X"00",X"73",X"30",X"BB",X"BD",X"C3",X"33",
		X"3E",X"00",X"0A",X"BA",X"C7",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"09",X"01",X"05",
		X"FF",X"FF",X"09",X"E7",X"FB",X"80",X"09",X"06",X"03",X"55",X"50",X"05",X"00",X"00",X"00",X"00",
		X"55",X"55",X"55",X"55",X"50",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"0A",X"01",X"0A",X"01",
		X"0A",X"01",X"0A",X"FF",X"FF",X"0A",X"0A",X"05",X"00",X"09",X"06",X"03",X"00",X"00",X"05",X"00",
		X"55",X"50",X"55",X"55",X"55",X"55",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"0A",X"00",X"0A",X"01",X"0A",X"FF",X"FF",X"0A",X"2D",X"FC",X"80",X"01",X"06",X"03",X"33",
		X"70",X"03",X"00",X"72",X"00",X"0E",X"33",X"33",X"19",X"29",X"E0",X"00",X"00",X"0E",X"D7",X"7E",
		X"00",X"00",X"09",X"01",X"0A",X"05",X"09",X"FF",X"FF",X"0A",X"4E",X"06",X"80",X"01",X"06",X"03",
		X"02",X"70",X"03",X"00",X"73",X"30",X"E9",X"29",X"13",X"33",X"3E",X"00",X"0E",X"77",X"DE",X"00",
		X"00",X"00",X"01",X"0A",X"00",X"09",X"01",X"05",X"FF",X"FF",X"0A",X"BA",X"FF",X"00",X"F9",X"0A",
		X"F6",X"00",X"80",X"F8",X"0B",X"24",X"04",X"00",X"F6",X"0B",X"52",X"07",X"80",X"FA",X"0B",X"80",
		X"0C",X"00",X"FD",X"0B",X"AE",X"07",X"80",X"01",X"0B",X"DC",X"04",X"00",X"05",X"0C",X"0A",X"00",
		X"80",X"01",X"0A",X"BA",X"02",X"00",X"F9",X"0C",X"0A",X"FE",X"00",X"FA",X"0B",X"DC",X"FA",X"80",
		X"F6",X"0B",X"AE",X"F7",X"00",X"FA",X"0B",X"80",X"F4",X"80",X"FD",X"0B",X"52",X"F7",X"00",X"01",
		X"0B",X"24",X"FA",X"80",X"04",X"0A",X"F6",X"FE",X"00",X"01",X"05",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"B5",X"75",X"B0",X"00",X"0C",X"9C",X"5C",X"4C",X"00",
		X"04",X"14",X"44",X"44",X"00",X"0C",X"4C",X"44",X"4C",X"00",X"0E",X"4C",X"4C",X"CE",X"00",X"00",
		X"EE",X"CE",X"E0",X"00",X"00",X"00",X"04",X"04",X"02",X"06",X"01",X"07",X"01",X"07",X"01",X"07",
		X"01",X"07",X"02",X"06",X"FF",X"FF",X"04",X"07",X"0E",X"4C",X"50",X"00",X"C1",X"9C",X"BE",X"50",
		X"44",X"C4",X"55",X"00",X"CE",X"44",X"CC",X"50",X"EC",X"44",X"47",X"C0",X"0C",X"CC",X"CC",X"E0",
		X"00",X"EE",X"CE",X"00",X"01",X"04",X"00",X"06",X"00",X"05",X"00",X"06",X"00",X"06",X"01",X"06",
		X"02",X"05",X"FF",X"FF",X"04",X"07",X"0E",X"C4",X"E0",X"00",X"E4",X"19",X"4B",X"00",X"CC",X"C4",
		X"E5",X"00",X"C4",X"44",X"5E",X"50",X"CC",X"44",X"E5",X"00",X"EC",X"4C",X"CB",X"00",X"0E",X"7C",
		X"E0",X"00",X"01",X"04",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"05",X"00",X"05",X"01",X"04",
		X"FF",X"FF",X"04",X"07",X"00",X"EC",X"CE",X"00",X"0C",X"C1",X"94",X"E0",X"E4",X"44",X"C4",X"C0",
		X"44",X"44",X"4C",X"E0",X"CC",X"4C",X"5B",X"50",X"EC",X"CE",X"5E",X"00",X"0E",X"C5",X"05",X"00",
		X"02",X"05",X"01",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"01",X"05",X"FF",X"FF",
		X"04",X"07",X"0E",X"4C",X"EE",X"00",X"C1",X"44",X"CC",X"C0",X"49",X"44",X"C4",X"C0",X"44",X"44",
		X"44",X"40",X"E7",X"C5",X"CC",X"E0",X"0B",X"5E",X"5B",X"00",X"00",X"05",X"00",X"00",X"01",X"05",
		X"00",X"06",X"00",X"06",X"00",X"06",X"00",X"06",X"01",X"05",X"03",X"03",X"FF",X"FF",X"04",X"07",
		X"0E",X"4C",X"E0",X"00",X"E9",X"14",X"CC",X"00",X"C4",X"44",X"4C",X"E0",X"EC",X"44",X"4E",X"C0",
		X"5B",X"5E",X"CC",X"C0",X"0E",X"5E",X"CC",X"E0",X"05",X"05",X"CE",X"00",X"01",X"04",X"00",X"05",
		X"00",X"06",X"00",X"06",X"00",X"06",X"01",X"06",X"01",X"05",X"FF",X"FF",X"04",X"07",X"00",X"C4",
		X"CC",X"00",X"0B",X"41",X"44",X"E0",X"05",X"C4",X"44",X"40",X"54",X"54",X"44",X"C0",X"05",X"E4",
		X"CC",X"E0",X"0B",X"C4",X"4C",X"E0",X"00",X"E7",X"CE",X"00",X"02",X"05",X"01",X"06",X"01",X"06",
		X"00",X"06",X"01",X"06",X"01",X"06",X"02",X"05",X"FF",X"FF",X"04",X"07",X"00",X"5C",X"4E",X"00",
		X"57",X"B1",X"94",X"C0",X"05",X"59",X"44",X"40",X"5E",X"44",X"44",X"C0",X"C4",X"C4",X"7C",X"E0",
		X"EC",X"CC",X"CC",X"00",X"0E",X"CC",X"E0",X"00",X"02",X"05",X"00",X"06",X"01",X"06",X"00",X"06",
		X"00",X"06",X"00",X"05",X"01",X"04",X"FF",X"FF",X"0C",X"60",X"FD",X"80",X"F9",X"0C",X"AC",X"00",
		X"80",X"FA",X"0C",X"F8",X"04",X"00",X"F6",X"0D",X"3E",X"07",X"80",X"FA",X"0D",X"8F",X"0C",X"00",
		X"FD",X"0D",X"CB",X"07",X"80",X"01",X"0E",X"17",X"04",X"00",X"05",X"0E",X"5D",X"00",X"80",X"01",
		X"07",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",
		X"00",X"00",X"00",X"86",X"80",X"00",X"00",X"06",X"80",X"0F",X"66",X"6D",X"00",X"00",X"00",X"86",
		X"81",X"66",X"11",X"10",X"00",X"00",X"06",X"66",X"81",X"90",X"12",X"00",X"00",X"88",X"F8",X"8D",
		X"11",X"19",X"00",X"08",X"F0",X"0F",X"88",X"11",X"B0",X"00",X"00",X"00",X"05",X"06",X"06",X"08",
		X"01",X"09",X"02",X"0A",X"03",X"0B",X"02",X"0B",X"01",X"0A",X"FF",X"FF",X"06",X"09",X"00",X"00",
		X"F6",X"D1",X"D2",X"00",X"00",X"06",X"66",X"10",X"11",X"90",X"00",X"6F",X"66",X"17",X"11",X"00",
		X"00",X"00",X"61",X"81",X"1B",X"00",X"60",X"00",X"66",X"88",X"80",X"00",X"06",X"66",X"68",X"88",
		X"00",X"00",X"00",X"F8",X"8F",X"F0",X"00",X"00",X"00",X"08",X"80",X"00",X"00",X"00",X"08",X"88",
		X"00",X"00",X"00",X"00",X"04",X"09",X"03",X"0A",X"02",X"09",X"04",X"09",X"00",X"08",X"01",X"07",
		X"02",X"06",X"03",X"04",X"01",X"03",X"FF",X"FF",X"04",X"0B",X"00",X"00",X"29",X"00",X"00",X"01",
		X"11",X"B0",X"00",X"D1",X"01",X"10",X"08",X"61",X"91",X"10",X"F6",X"16",X"1D",X"80",X"88",X"66",
		X"88",X"80",X"80",X"F6",X"88",X"F0",X"00",X"06",X"6F",X"00",X"00",X"06",X"88",X"00",X"00",X"88",
		X"08",X"F0",X"00",X"60",X"00",X"80",X"04",X"05",X"03",X"06",X"02",X"06",X"01",X"06",X"00",X"06",
		X"00",X"06",X"00",X"06",X"03",X"05",X"03",X"05",X"02",X"06",X"02",X"06",X"FF",X"FF",X"05",X"0B",
		X"09",X"00",X"00",X"00",X"00",X"21",X"1D",X"00",X"00",X"00",X"D1",X"11",X"6F",X"00",X"00",X"10",
		X"91",X"66",X"00",X"00",X"D1",X"16",X"66",X"F0",X"00",X"68",X"81",X"66",X"60",X"00",X"F8",X"88",
		X"86",X"68",X"00",X"08",X"F0",X"08",X"88",X"F0",X"00",X"60",X"06",X"F0",X"80",X"00",X"00",X"08",
		X"00",X"80",X"00",X"00",X"80",X"00",X"00",X"01",X"01",X"00",X"03",X"00",X"05",X"00",X"05",X"00",
		X"06",X"00",X"06",X"00",X"07",X"01",X"08",X"02",X"08",X"05",X"08",X"04",X"04",X"FF",X"FF",X"06",
		X"07",X"0B",X"11",X"D6",X"80",X"08",X"60",X"21",X"11",X"16",X"66",X"68",X"00",X"91",X"09",X"18",
		X"16",X"80",X"00",X"01",X"11",X"88",X"88",X"88",X"00",X"00",X"D8",X"88",X"F0",X"0F",X"80",X"00",
		X"0F",X"88",X"00",X"00",X"00",X"00",X"00",X"0F",X"80",X"00",X"00",X"01",X"0A",X"00",X"09",X"00",
		X"08",X"01",X"09",X"02",X"0A",X"03",X"05",X"05",X"06",X"FF",X"FF",X"06",X"09",X"00",X"00",X"00",
		X"08",X"66",X"00",X"00",X"00",X"00",X"68",X"00",X"00",X"00",X"00",X"86",X"66",X"F0",X"00",X"00",
		X"06",X"16",X"F8",X"88",X"00",X"00",X"66",X"68",X"80",X"00",X"80",X"0D",X"11",X"88",X"80",X"00",
		X"00",X"01",X"19",X"18",X"8F",X"80",X"00",X"21",X"10",X"18",X"88",X"00",X"00",X"02",X"D1",X"D8",
		X"F0",X"00",X"00",X"07",X"09",X"06",X"07",X"04",X"08",X"03",X"09",X"02",X"0A",X"01",X"06",X"01",
		X"08",X"00",X"07",X"01",X"06",X"FF",X"FF",X"04",X"0B",X"60",X"00",X"60",X"00",X"88",X"08",X"F0",
		X"00",X"06",X"88",X"00",X"00",X"06",X"68",X"00",X"00",X"F1",X"66",X"F0",X"80",X"66",X"86",X"88",
		X"80",X"61",X"D8",X"88",X"00",X"11",X"91",X"88",X"00",X"11",X"01",X"D0",X"00",X"B1",X"11",X"00",
		X"00",X"02",X"90",X"00",X"00",X"00",X"04",X"00",X"04",X"01",X"03",X"01",X"03",X"00",X"06",X"00",
		X"06",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"03",X"01",X"02",X"FF",X"FF",X"05",X"0B",X"00",
		X"00",X"60",X"00",X"00",X"60",X"06",X"00",X"00",X"00",X"60",X"F8",X"00",X"60",X"00",X"86",X"86",
		X"00",X"F6",X"00",X"06",X"66",X"66",X"66",X"F0",X"00",X"86",X"16",X"88",X"80",X"00",X"88",X"88",
		X"11",X"D0",X"00",X"08",X"81",X"20",X"10",X"00",X"0F",X"81",X"11",X"10",X"00",X"00",X"FD",X"11",
		X"20",X"00",X"00",X"00",X"02",X"00",X"04",X"04",X"00",X"03",X"00",X"06",X"00",X"07",X"01",X"08",
		X"02",X"08",X"02",X"08",X"03",X"08",X"03",X"08",X"04",X"08",X"07",X"07",X"FF",X"FF",X"0E",X"D6",
		X"01",X"80",X"F9",X"10",X"D3",X"FE",X"00",X"FA",X"10",X"8D",X"FA",X"80",X"F6",X"10",X"41",X"F7",
		X"00",X"FA",X"10",X"05",X"F4",X"80",X"FD",X"0F",X"B4",X"F7",X"00",X"01",X"0F",X"6E",X"FA",X"80",
		X"04",X"0F",X"22",X"FE",X"00",X"01",X"07",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"86",X"00",X"00",X"00",X"00",X"00",X"86",X"80",X"00",X"00",X"00",X"00",X"0D",X"61",
		X"6F",X"00",X"86",X"00",X"00",X"D1",X"16",X"66",X"86",X"80",X"00",X"02",X"10",X"91",X"88",X"66",
		X"00",X"00",X"09",X"11",X"1D",X"88",X"F8",X"80",X"00",X"00",X"B1",X"18",X"8F",X"00",X"F8",X"00",
		X"00",X"00",X"06",X"07",X"04",X"06",X"03",X"0B",X"02",X"0A",X"01",X"09",X"01",X"0A",X"02",X"0B",
		X"FF",X"FF",X"06",X"09",X"02",X"D1",X"D6",X"F0",X"00",X"00",X"21",X"10",X"16",X"68",X"00",X"00",
		X"01",X"19",X"16",X"66",X"60",X"00",X"0B",X"11",X"81",X"60",X"00",X"00",X"00",X"88",X"86",X"60",
		X"00",X"60",X"00",X"08",X"88",X"66",X"66",X"00",X"00",X"00",X"F8",X"88",X"80",X"00",X"00",X"00",
		X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"0F",X"88",X"00",X"01",X"06",X"00",X"07",X"01",X"08",
		X"01",X"06",X"02",X"0A",X"03",X"09",X"04",X"08",X"06",X"07",X"07",X"09",X"FF",X"FF",X"04",X"0B",
		X"02",X"90",X"00",X"00",X"B1",X"11",X"00",X"00",X"11",X"01",X"D0",X"00",X"11",X"91",X"8F",X"00",
		X"61",X"18",X"86",X"00",X"66",X"86",X"88",X"80",X"F6",X"68",X"F0",X"80",X"08",X"6F",X"00",X"00",
		X"08",X"68",X"00",X"00",X"86",X"08",X"F0",X"00",X"60",X"00",X"60",X"00",X"01",X"02",X"00",X"03",
		X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"06",X"00",X"06",X"01",X"03",X"01",X"03",X"00",X"04",
		X"00",X"04",X"FF",X"FF",X"05",X"0B",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"0D",X"11",X"20",
		X"00",X"00",X"61",X"11",X"10",X"00",X"06",X"61",X"10",X"10",X"00",X"F1",X"68",X"17",X"D0",X"00",
		X"66",X"68",X"68",X"80",X"08",X"68",X"88",X"88",X"F0",X"86",X"88",X"00",X"8F",X"00",X"60",X"88",
		X"00",X"80",X"00",X"60",X"06",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"07",X"07",X"05",
		X"08",X"04",X"08",X"03",X"08",X"02",X"08",X"02",X"08",X"01",X"08",X"00",X"07",X"00",X"06",X"00",
		X"03",X"04",X"04",X"FF",X"FF",X"06",X"07",X"68",X"00",X"F6",X"6D",X"1B",X"00",X"08",X"88",X"66",
		X"11",X"11",X"90",X"00",X"66",X"16",X"19",X"01",X"20",X"08",X"88",X"88",X"81",X"11",X"00",X"6F",
		X"00",X"F8",X"88",X"D0",X"00",X"00",X"00",X"08",X"8F",X"00",X"00",X"00",X"00",X"88",X"00",X"00",
		X"00",X"00",X"09",X"01",X"0A",X"02",X"0A",X"01",X"09",X"00",X"08",X"05",X"07",X"04",X"05",X"FF",
		X"FF",X"06",X"09",X"06",X"8F",X"00",X"00",X"00",X"00",X"00",X"06",X"80",X"00",X"00",X"00",X"00",
		X"F8",X"66",X"80",X"00",X"00",X"06",X"68",X"66",X"66",X"00",X"00",X"60",X"00",X"F1",X"66",X"80",
		X"00",X"00",X"00",X"86",X"81",X"1B",X"00",X"00",X"68",X"88",X"12",X"11",X"00",X"00",X"08",X"88",
		X"70",X"11",X"20",X"00",X"00",X"F8",X"D1",X"D2",X"00",X"01",X"03",X"03",X"04",X"02",X"06",X"01",
		X"07",X"00",X"08",X"04",X"09",X"02",X"09",X"03",X"0A",X"04",X"09",X"FF",X"FF",X"04",X"0B",X"00",
		X"60",X"00",X"60",X"00",X"88",X"08",X"F0",X"00",X"06",X"68",X"00",X"00",X"06",X"88",X"00",X"60",
		X"86",X"68",X"F0",X"86",X"16",X"88",X"80",X"06",X"88",X"1D",X"60",X"0F",X"81",X"91",X"D0",X"00",
		X"D1",X"01",X"10",X"00",X"01",X"11",X"D0",X"00",X"00",X"29",X"00",X"02",X"06",X"02",X"06",X"03",
		X"05",X"03",X"05",X"00",X"06",X"00",X"06",X"01",X"06",X"01",X"06",X"02",X"06",X"03",X"06",X"04",
		X"05",X"FF",X"FF",X"05",X"0B",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"06",X"00",X"60",X"00",
		X"60",X"06",X"80",X"80",X"08",X"60",X"08",X"88",X"F0",X"F6",X"66",X"86",X"88",X"00",X"66",X"66",
		X"18",X"80",X"00",X"D1",X"18",X"88",X"F0",X"00",X"10",X"71",X"88",X"00",X"00",X"D1",X"11",X"80",
		X"00",X"00",X"21",X"1B",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"04",X"04",X"05",X"08",
		X"02",X"08",X"01",X"08",X"00",X"07",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"04",X"00",X"03",
		X"01",X"01",X"FF",X"FF",X"11",X"74",X"FD",X"00",X"FA",X"11",X"BE",X"00",X"80",X"F8",X"12",X"0A",
		X"04",X"00",X"F6",X"12",X"56",X"07",X"80",X"FA",X"12",X"A0",X"0C",X"00",X"FD",X"12",X"DA",X"07",
		X"80",X"01",X"13",X"24",X"04",X"00",X"05",X"13",X"70",X"00",X"80",X"01",X"11",X"74",X"01",X"80",
		X"FA",X"13",X"70",X"FE",X"00",X"FA",X"13",X"24",X"FA",X"80",X"F6",X"12",X"DA",X"F7",X"00",X"FA",
		X"12",X"A0",X"F4",X"80",X"FD",X"12",X"56",X"F7",X"00",X"01",X"12",X"0A",X"FA",X"80",X"04",X"11",
		X"BE",X"FE",X"00",X"01",X"08",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"21",X"21",X"00",X"00",X"00",X"00",X"12",
		X"11",X"12",X"12",X"21",X"00",X"00",X"01",X"11",X"21",X"9D",X"19",X"72",X"10",X"00",X"0D",X"CC",
		X"19",X"EC",X"21",X"CC",X"D0",X"00",X"00",X"0E",X"CC",X"CC",X"CC",X"E0",X"00",X"00",X"00",X"00",
		X"06",X"07",X"04",X"09",X"02",X"0B",X"01",X"0C",X"01",X"0C",X"03",X"0A",X"FF",X"FF",X"06",X"09",
		X"11",X"19",X"00",X"00",X"00",X"00",X"04",X"D1",X"11",X"04",X"00",X"00",X"0C",X"E2",X"11",X"1C",
		X"00",X"00",X"00",X"C1",X"9D",X"11",X"00",X"00",X"00",X"02",X"E7",X"12",X"B0",X"00",X"00",X"00",
		X"CC",X"1D",X"20",X"00",X"00",X"00",X"0C",X"17",X"10",X"00",X"00",X"00",X"00",X"EC",X"1D",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"03",X"01",X"07",X"01",X"07",X"02",X"07",X"03",X"08",
		X"04",X"08",X"05",X"08",X"06",X"09",X"08",X"08",X"FF",X"FF",X"04",X"0C",X"0D",X"10",X"00",X"00",
		X"0C",X"11",X"00",X"00",X"CE",X"12",X"00",X"00",X"C1",X"21",X"10",X"00",X"49",X"11",X"10",X"00",
		X"4E",X"D1",X"14",X"00",X"CC",X"92",X"7C",X"00",X"C2",X"1D",X"20",X"00",X"C1",X"D1",X"10",X"00",
		X"EC",X"72",X"00",X"00",X"0E",X"D1",X"00",X"00",X"0D",X"10",X"00",X"00",X"01",X"02",X"01",X"03",
		X"00",X"03",X"00",X"04",X"00",X"04",X"00",X"05",X"00",X"05",X"00",X"04",X"00",X"04",X"00",X"03",
		X"01",X"03",X"01",X"02",X"FF",X"FF",X"05",X"0A",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",
		X"CC",X"70",X"00",X"00",X"0C",X"EB",X"10",X"00",X"00",X"21",X"91",X"90",X"00",X"0C",X"E9",X"11",
		X"00",X"00",X"CC",X"D1",X"11",X"00",X"0E",X"11",X"1D",X"10",X"00",X"0C",X"7D",X"21",X"04",X"00",
		X"19",X"12",X"B0",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"08",X"08",X"06",X"08",X"05",X"08",
		X"04",X"08",X"03",X"07",X"02",X"07",X"01",X"06",X"01",X"07",X"00",X"04",X"01",X"01",X"FF",X"FF",
		X"07",X"06",X"00",X"EC",X"44",X"CC",X"CC",X"00",X"00",X"DC",X"C1",X"2E",X"C9",X"1E",X"CD",X"00",
		X"11",X"12",X"1D",X"71",X"D7",X"21",X"00",X"01",X"21",X"11",X"21",X"91",X"10",X"00",X"00",X"01",
		X"91",X"12",X"10",X"00",X"00",X"00",X"00",X"04",X"C0",X"00",X"00",X"00",X"02",X"09",X"00",X"0B",
		X"00",X"0B",X"01",X"0A",X"03",X"08",X"05",X"06",X"FF",X"FF",X"05",X"0A",X"10",X"00",X"00",X"00",
		X"00",X"1C",X"C0",X"00",X"00",X"00",X"DD",X"EC",X"00",X"00",X"00",X"11",X"91",X"20",X"00",X"00",
		X"E1",X"1D",X"EC",X"00",X"00",X"01",X"12",X"DC",X"C0",X"00",X"04",X"12",X"11",X"1E",X"00",X"00",
		X"01",X"2D",X"EC",X"00",X"00",X"00",X"B2",X"11",X"D0",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",
		X"00",X"02",X"00",X"03",X"00",X"04",X"00",X"05",X"01",X"06",X"01",X"07",X"03",X"07",X"04",X"08",
		X"07",X"07",X"FF",X"FF",X"04",X"0C",X"00",X"01",X"D0",X"00",X"00",X"11",X"C0",X"00",X"00",X"11",
		X"EC",X"00",X"09",X"12",X"1C",X"00",X"01",X"11",X"2C",X"00",X"42",X"1D",X"CC",X"00",X"C1",X"29",
		X"EC",X"00",X"02",X"D1",X"1C",X"00",X"01",X"2D",X"2C",X"00",X"00",X"17",X"CE",X"00",X"00",X"1D",
		X"E0",X"00",X"00",X"01",X"D0",X"00",X"03",X"04",X"02",X"04",X"02",X"05",X"01",X"05",X"01",X"05",
		X"00",X"05",X"00",X"05",X"01",X"05",X"01",X"05",X"02",X"05",X"02",X"04",X"03",X"04",X"FF",X"FF",
		X"06",X"09",X"00",X"00",X"07",X"11",X"DD",X"00",X"00",X"40",X"11",X"1D",X"C0",X"00",X"00",X"C1",
		X"11",X"2E",X"C0",X"00",X"00",X"1D",X"71",X"1C",X"00",X"00",X"0B",X"21",X"9E",X"20",X"00",X"00",
		X"01",X"D1",X"CC",X"00",X"00",X"00",X"0D",X"71",X"C0",X"00",X"00",X"00",X"B1",X"CE",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"05",X"09",X"02",X"08",X"02",X"08",X"02",X"07",
		X"01",X"06",X"01",X"05",X"01",X"04",X"00",X"03",X"01",X"01",X"FF",X"FF",X"14",X"0C",X"FE",X"80",
		X"FC",X"14",X"38",X"00",X"80",X"F9",X"14",X"7B",X"04",X"00",X"F6",X"14",X"AC",X"07",X"80",X"FA",
		X"14",X"EF",X"0C",X"00",X"FD",X"15",X"0F",X"07",X"80",X"01",X"15",X"52",X"04",X"00",X"05",X"15",
		X"83",X"00",X"80",X"01",X"14",X"0C",X"01",X"80",X"FC",X"15",X"83",X"FE",X"00",X"FA",X"15",X"52",
		X"FA",X"80",X"F6",X"15",X"0F",X"F7",X"00",X"FA",X"14",X"EF",X"F4",X"80",X"FD",X"14",X"AC",X"F7",
		X"00",X"01",X"14",X"7B",X"FA",X"80",X"04",X"14",X"38",X"FE",X"00",X"01",X"06",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"02",X"00",X"01",X"97",X"00",X"0E",X"92",X"00",
		X"07",X"22",X"22",X"22",X"27",X"00",X"00",X"E7",X"22",X"27",X"E0",X"00",X"00",X"00",X"01",X"09",
		X"01",X"09",X"01",X"09",X"02",X"08",X"FF",X"FF",X"05",X"09",X"02",X"00",X"00",X"00",X"00",X"79",
		X"00",X"00",X"00",X"00",X"12",X"70",X"00",X"00",X"00",X"72",X"90",X"00",X"00",X"00",X"E2",X"77",
		X"00",X"00",X"00",X"07",X"22",X"70",X"00",X"00",X"00",X"79",X"29",X"E0",X"00",X"00",X"07",X"97",
		X"99",X"90",X"00",X"00",X"E7",X"97",X"00",X"01",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"00",
		X"03",X"01",X"04",X"02",X"06",X"03",X"08",X"04",X"07",X"FF",X"FF",X"03",X"09",X"07",X"22",X"00",
		X"E1",X"20",X"00",X"72",X"E0",X"00",X"22",X"00",X"00",X"22",X"00",X"00",X"22",X"00",X"00",X"79",
		X"70",X"00",X"E9",X"20",X"00",X"0E",X"92",X"00",X"01",X"03",X"00",X"02",X"00",X"02",X"00",X"01",
		X"00",X"01",X"00",X"01",X"00",X"02",X"00",X"02",X"01",X"03",X"FF",X"FF",X"05",X"09",X"00",X"00",
		X"07",X"97",X"00",X"00",X"07",X"21",X"22",X"90",X"00",X"72",X"27",X"E0",X"00",X"07",X"22",X"70",
		X"00",X"00",X"E2",X"27",X"00",X"00",X"00",X"77",X"90",X"00",X"00",X"00",X"92",X"E0",X"00",X"00",
		X"00",X"79",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"05",X"07",X"03",X"08",X"02",
		X"06",X"01",X"04",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"01",X"01",X"01",X"FF",X"FF",X"05",
		X"04",X"0E",X"72",X"22",X"7E",X"00",X"71",X"22",X"22",X"22",X"70",X"29",X"E0",X"00",X"E9",X"90",
		X"20",X"00",X"00",X"00",X"20",X"01",X"07",X"00",X"08",X"00",X"08",X"00",X"08",X"FF",X"FF",X"05",
		X"09",X"07",X"97",X"00",X"00",X"00",X"92",X"12",X"27",X"00",X"00",X"00",X"E9",X"72",X"70",X"00",
		X"00",X"00",X"79",X"27",X"00",X"00",X"00",X"07",X"22",X"E0",X"00",X"00",X"00",X"77",X"70",X"00",
		X"00",X"00",X"E9",X"90",X"00",X"00",X"00",X"09",X"70",X"00",X"00",X"00",X"02",X"00",X"01",X"03",
		X"00",X"05",X"02",X"06",X"04",X"07",X"05",X"08",X"06",X"08",X"06",X"08",X"07",X"08",X"07",X"07",
		X"FF",X"FF",X"03",X"09",X"22",X"70",X"00",X"02",X"1E",X"00",X"0E",X"27",X"00",X"00",X"22",X"00",
		X"00",X"22",X"00",X"00",X"92",X"00",X"07",X"27",X"00",X"02",X"9E",X"00",X"29",X"E0",X"00",X"00",
		X"02",X"01",X"03",X"01",X"03",X"02",X"03",X"02",X"03",X"02",X"03",X"01",X"03",X"01",X"03",X"00",
		X"02",X"FF",X"FF",X"05",X"09",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"02",X"E0",X"00",
		X"00",X"00",X"71",X"90",X"00",X"00",X"00",X"22",X"70",X"00",X"00",X"07",X"79",X"E0",X"00",X"00",
		X"72",X"97",X"00",X"00",X"E9",X"29",X"70",X"00",X"22",X"27",X"97",X"00",X"00",X"07",X"97",X"E0",
		X"00",X"00",X"07",X"07",X"07",X"08",X"06",X"08",X"06",X"08",X"05",X"08",X"04",X"07",X"02",X"06",
		X"00",X"05",X"01",X"04",X"FF",X"FF",X"16",X"16",X"FF",X"80",X"F9",X"16",X"52",X"00",X"80",X"F7",
		X"16",X"7A",X"04",X"00",X"F7",X"16",X"A2",X"07",X"80",X"F7",X"16",X"CA",X"0C",X"00",X"F8",X"16",
		X"F8",X"07",X"80",X"01",X"17",X"20",X"04",X"00",X"05",X"17",X"48",X"00",X"80",X"01",X"16",X"16",
		X"02",X"00",X"F9",X"17",X"48",X"FE",X"00",X"FA",X"17",X"20",X"FA",X"80",X"F6",X"16",X"F8",X"F7",
		X"00",X"FA",X"16",X"CA",X"F4",X"80",X"FD",X"16",X"A2",X"F7",X"00",X"01",X"16",X"7A",X"FA",X"80",
		X"04",X"16",X"52",X"FE",X"00",X"01",X"05",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"10",
		X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"0B",X"11",X"11",X"B0",X"00",X"0D",X"11",X"11",X"D0",
		X"00",X"0D",X"11",X"1D",X"D0",X"00",X"0B",X"11",X"DD",X"A0",X"00",X"00",X"B1",X"DB",X"00",X"00",
		X"00",X"00",X"03",X"04",X"02",X"05",X"01",X"06",X"01",X"06",X"01",X"06",X"01",X"06",X"02",X"05",
		X"FF",X"FF",X"04",X"06",X"00",X"BD",X"11",X"D0",X"01",X"11",X"11",X"10",X"D1",X"11",X"11",X"D0",
		X"DD",X"11",X"11",X"B0",X"BD",X"D1",X"1D",X"00",X"0B",X"DD",X"B0",X"00",X"02",X"06",X"01",X"06",
		X"00",X"06",X"00",X"06",X"00",X"05",X"01",X"04",X"FF",X"FF",X"04",X"06",X"0B",X"DD",X"B0",X"00",
		X"B1",X"11",X"11",X"00",X"11",X"11",X"11",X"10",X"D1",X"11",X"11",X"10",X"BD",X"D1",X"11",X"00",
		X"0A",X"DD",X"B0",X"00",X"01",X"04",X"00",X"05",X"00",X"06",X"00",X"06",X"00",X"05",X"01",X"04",
		X"FF",X"FF",X"04",X"06",X"0B",X"DD",X"B0",X"00",X"BD",X"11",X"1D",X"00",X"D1",X"11",X"11",X"B0",
		X"BD",X"11",X"11",X"D0",X"0D",X"D1",X"11",X"10",X"00",X"BD",X"11",X"D0",X"01",X"04",X"00",X"05",
		X"00",X"06",X"00",X"06",X"01",X"06",X"02",X"06",X"FF",X"FF",X"04",X"07",X"0B",X"1D",X"B0",X"00",
		X"B1",X"1D",X"DA",X"00",X"D1",X"11",X"DD",X"00",X"D1",X"11",X"1D",X"00",X"B1",X"11",X"1B",X"00",
		X"01",X"11",X"10",X"00",X"00",X"11",X"00",X"00",X"01",X"04",X"00",X"05",X"00",X"05",X"00",X"05",
		X"00",X"05",X"01",X"04",X"02",X"03",X"FF",X"FF",X"04",X"06",X"00",X"BD",X"DB",X"00",X"0D",X"11",
		X"1D",X"B0",X"B1",X"11",X"1D",X"D0",X"D1",X"11",X"1D",X"B0",X"11",X"11",X"DD",X"00",X"D1",X"1D",
		X"B0",X"00",X"02",X"05",X"01",X"06",X"00",X"06",X"00",X"06",X"00",X"05",X"00",X"04",X"FF",X"FF",
		X"04",X"06",X"00",X"BD",X"DB",X"00",X"01",X"11",X"11",X"B0",X"11",X"11",X"11",X"D0",X"11",X"11",
		X"1D",X"D0",X"01",X"11",X"DD",X"A0",X"00",X"BD",X"DA",X"00",X"02",X"05",X"01",X"06",X"00",X"06",
		X"00",X"06",X"01",X"06",X"02",X"05",X"FF",X"FF",X"04",X"06",X"D1",X"1D",X"B0",X"00",X"11",X"11",
		X"1D",X"00",X"D1",X"11",X"11",X"D0",X"B1",X"11",X"1D",X"D0",X"0D",X"11",X"1D",X"B0",X"00",X"BD",
		X"DB",X"00",X"00",X"04",X"00",X"05",X"00",X"06",X"00",X"06",X"01",X"06",X"02",X"05",X"FF",X"FF",
		X"17",X"C0",X"02",X"80",X"FC",X"17",X"C0",X"FE",X"00",X"FA",X"17",X"C0",X"FA",X"80",X"F6",X"17",
		X"C0",X"F7",X"00",X"FA",X"17",X"C0",X"F4",X"80",X"FD",X"17",X"C0",X"F7",X"00",X"01",X"17",X"C0",
		X"FA",X"80",X"04",X"17",X"C0",X"FE",X"00",X"01",X"17",X"C0",X"00",X"00",X"FC",X"17",X"C0",X"00",
		X"80",X"FA",X"17",X"C0",X"04",X"00",X"F6",X"17",X"C0",X"07",X"80",X"FA",X"17",X"C0",X"0C",X"00",
		X"FD",X"17",X"C0",X"07",X"80",X"01",X"17",X"C0",X"04",X"00",X"05",X"17",X"C0",X"00",X"80",X"01",
		X"04",X"05",X"00",X"D1",X"00",X"00",X"00",X"11",X"D0",X"00",X"10",X"17",X"91",X"B0",X"11",X"19",
		X"91",X"10",X"01",X"10",X"01",X"00",X"02",X"03",X"02",X"04",X"00",X"06",X"00",X"06",X"01",X"05",
		X"FF",X"FF",X"19",X"1D",X"2A",X"76",X"22",X"83",X"AA",X"3B",X"CD",X"93",X"F5",X"D5",X"1D",X"88",
		X"A0",X"D7",X"71",X"DE",X"6F",X"E4",X"AF",X"EB",X"B8",X"EF",X"22",X"28",X"3A",X"D3",X"7A",X"EB",
		X"0E",X"B4",X"DE",X"B7",X"11",X"41",X"CD",X"F7",X"69",X"77",X"AE",X"A0",X"EF",X"37",X"DD",X"A5",
		X"DE",X"A2",X"28",X"37",X"D4",X"6B",X"76",X"AB",X"9B",X"EA",X"35",X"BB",X"89",X"A3",X"5B",X"61",
		X"C2",X"AE",X"90",X"70",X"AB",X"A6",X"1A",X"DC",X"5C",X"34",X"C2",X"44",X"58",X"1C",X"98",X"48",
		X"8A",X"2E",X"38",X"AB",X"1B",X"EE",X"F5",X"8E",X"0D",X"3E",X"63",X"49",X"75",X"17",X"1C",X"D7",
		X"75",X"8D",X"F5",X"A6",X"FA",X"43",X"2A",X"90",X"FB",X"B6",X"9D",X"D4",X"5C",X"73",X"5D",X"D6",
		X"37",X"DE",X"6F",X"5C",X"21",X"F7",X"49",X"98",X"A6",X"D7",X"48",X"7C",X"D6",X"F9",X"DD",X"45",
		X"C7",X"35",X"D4",X"4B",X"37",X"AE",X"3B",X"EF",X"8C",X"3E",X"EB",X"BE",X"6B",X"7C",X"EE",X"A2",
		X"E3",X"9A",X"7B",X"CD",X"EB",X"8C",X"FA",X"20",X"7A",X"CF",X"9A",X"DF",X"3B",X"A8",X"B8",X"44",
		X"F7",X"9B",X"D7",X"15",X"F4",X"48",X"F5",X"5F",X"35",X"BE",X"6F",X"51",X"20",X"10",X"B9",X"BD",
		X"71",X"1F",X"7C",X"24",X"7D",X"D4",X"7C",X"D6",X"DA",X"76",X"26",X"0D",X"F7",X"9B",X"D7",X"11",
		X"E8",X"50",X"E9",X"1F",X"35",X"BE",X"2D",X"E7",X"62",X"60",X"DF",X"79",X"BD",X"73",X"7D",X"F0",
		X"A1",X"F7",X"77",X"CD",X"6F",X"88",X"92",X"F2",X"25",X"0E",X"A4",X"D7",X"37",X"AE",X"6F",X"BE",
		X"14",X"3E",X"EE",X"F9",X"AD",X"F1",X"1E",X"BB",X"C8",X"92",X"3B",X"C5",X"BC",X"DE",X"B9",X"BE",
		X"8B",X"1E",X"EF",X"9A",X"DF",X"37",X"DD",X"77",X"91",X"24",X"73",X"BB",X"45",X"CD",X"EB",X"9B",
		X"E8",X"B1",X"EE",X"F9",X"AD",X"F3",X"7D",X"D7",X"79",X"12",X"47",X"3B",X"AE",X"EF",X"9B",X"D7",
		X"37",X"D1",X"63",X"DD",X"F3",X"5B",X"E6",X"FB",X"AE",X"F2",X"24",X"8E",X"77",X"5D",X"DF",X"37",
		X"AE",X"6F",X"A2",X"C7",X"BB",X"E6",X"B7",X"CD",X"F7",X"5D",X"E4",X"49",X"1C",X"EE",X"BB",X"BE",
		X"6F",X"5C",X"DF",X"7C",X"28",X"7D",X"DD",X"F3",X"5B",X"E6",X"FB",X"AE",X"F2",X"3C",X"DB",X"8E",
		X"77",X"5D",X"DF",X"37",X"AE",X"6F",X"BE",X"14",X"3E",X"EE",X"F9",X"AD",X"F3",X"7D",X"D7",X"78",
		X"E3",X"7C",X"8F",X"33",X"B6",X"1C",X"EE",X"BB",X"BE",X"6F",X"5C",X"47",X"A1",X"43",X"A4",X"7C",
		X"D6",X"F9",X"BE",X"EB",X"BC",X"61",X"BC",X"F2",X"3E",X"D6",X"5E",X"22",X"59",X"BD",X"71",X"1F",
		X"7C",X"24",X"7D",X"D4",X"7C",X"D6",X"F8",X"AB",X"A4",X"6D",X"7A",X"3E",X"D6",X"4B",X"5C",X"DE",
		X"B8",X"AF",X"A2",X"47",X"AA",X"F9",X"AD",X"A4",X"6A",X"CB",X"DA",X"F4",X"7D",X"AE",X"69",X"E6",
		X"B9",X"AE",X"6F",X"5C",X"67",X"D1",X"03",X"D6",X"7C",X"D6",X"F9",X"BE",X"74",X"87",X"ED",X"7A",
		X"3E",X"D7",X"34",X"B1",X"D7",X"37",X"AE",X"3B",X"EF",X"8C",X"3E",X"EB",X"BE",X"6B",X"69",X"37",
		X"C5",X"A8",X"FB",X"ED",X"7A",X"3E",X"D7",X"08",X"4B",X"79",X"BD",X"70",X"87",X"DD",X"26",X"62",
		X"9B",X"5D",X"21",X"F3",X"5B",X"E7",X"79",X"BE",X"3D",X"E6",X"BD",X"1F",X"6B",X"9A",X"66",X"D5",
		X"26",X"B9",X"BE",X"90",X"CA",X"A4",X"3E",X"EF",X"9A",X"32",X"77",X"DD",X"F4",X"7D",X"AE",X"75",
		X"DF",X"76",X"D7",X"83",X"4F",X"87",X"5D",X"F7",X"D1",X"F7",X"79",X"D4",X"44",X"D5",X"83",X"4B",
		X"87",X"5F",X"77",X"D1",X"F7",X"76",X"65",X"E6",X"B9",X"BE",X"EF",X"42",X"57",X"5B",X"EE",X"D6",
		X"19",X"77",X"DF",X"47",X"DD",X"E7",X"55",X"B5",X"59",X"BE",X"2B",X"D7",X"76",X"F5",X"1B",X"DD",
		X"F7",X"4A",X"F9",X"B3",X"27",X"77",X"DF",X"47",X"DD",X"DF",X"76",X"45",X"E6",X"F9",X"BE",X"2B",
		X"D2",X"D5",X"2D",X"54",X"AD",X"D2",X"BE",X"77",X"85",X"BE",X"EF",X"BE",X"8F",X"BB",X"B2",X"AA",
		X"CD",X"F1",X"5E",X"92",X"B9",X"4A",X"E5",X"2E",X"95",X"F3",X"BC",X"2D",X"F7",X"7D",X"F4",X"7D",
		X"DD",X"F7",X"65",X"5E",X"77",X"9B",X"EE",X"F4",X"95",X"0F",X"50",X"A5",X"43",X"D4",X"29",X"75",
		X"BE",X"EF",X"9A",X"E1",X"97",X"7D",X"F4",X"7D",X"DD",X"99",X"51",X"71",X"5E",X"92",X"E5",X"5E",
		X"52",X"E5",X"5E",X"52",X"B3",X"E1",X"D7",X"7D",X"F4",X"7D",X"DD",X"9F",X"78",X"AF",X"49",X"55",
		X"B5",X"56",X"97",X"4A",X"F8",X"7D",X"DF",X"7D",X"1F",X"23",X"10",X"5C",X"57",X"A7",X"BC",X"22",
		X"E9",X"5F",X"04",X"12",X"3F",X"47",X"DB",X"11",X"1D",X"CA",X"BD",X"77",X"5C",X"D7",X"35",X"CD",
		X"73",X"BA",X"57",X"9E",X"88",X"8D",X"FA",X"30",X"04",X"06",X"41",X"09",X"02",X"00",X"FD",X"DD",
		X"DF",X"0F",X"DB",X"FF",X"F8",X"FD",X"BF",X"FF",X"FF",X"D8",X"88",X"88",X"FF",X"08",X"B0",X"00",
		X"8F",X"08",X"B0",X"00",X"0D",X"04",X"06",X"41",X"09",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"D8",X"00",X"0D",X"BF",X"FF",X"00",X"DB",X"FF",X"FF",X"0D",X"BF",X"F8",X"8F",X"D8",X"88",
		X"80",X"0D",X"04",X"06",X"4F",X"09",X"02",X"00",X"00",X"00",X"00",X"DD",X"DD",X"F0",X"00",X"BF",
		X"FF",X"8F",X"00",X"FF",X"FF",X"F8",X"F0",X"F8",X"8F",X"FF",X"8F",X"80",X"08",X"88",X"88",X"04",
		X"06",X"4F",X"09",X"02",X"FD",X"DD",X"DF",X"00",X"DB",X"FF",X"F8",X"F0",X"BF",X"FF",X"FF",X"8F",
		X"FF",X"88",X"88",X"88",X"F8",X"00",X"08",X"B0",X"80",X"00",X"08",X"B0",X"02",X"03",X"40",X"2B",
		X"0A",X"FF",X"FB",X"FF",X"FB",X"FF",X"FB",X"02",X"03",X"40",X"2B",X"0A",X"DD",X"DD",X"DB",X"BB",
		X"DD",X"DD",X"04",X"08",X"52",X"27",X"0A",X"FF",X"DB",X"DF",X"FB",X"FF",X"FD",X"BD",X"FF",X"FF",
		X"FB",X"DB",X"DF",X"FF",X"FD",X"BB",X"BB",X"DD",X"6B",X"BD",X"BB",X"BB",X"BB",X"4F",X"BB",X"BB",
		X"DB",X"BB",X"BB",X"FF",X"FB",X"BB",X"BF",X"04",X"08",X"52",X"27",X"0A",X"FD",X"BD",X"FF",X"FB",
		X"FD",X"BD",X"FF",X"FF",X"FD",X"BD",X"FF",X"FF",X"BD",X"BB",X"BF",X"FF",X"DB",X"B6",X"BB",X"FF",
		X"BB",X"4F",X"BB",X"FF",X"DB",X"BB",X"BB",X"FF",X"FB",X"BB",X"BF",X"FF",X"04",X"02",X"48",X"31",
		X"0A",X"FF",X"F4",X"9F",X"FF",X"24",X"24",X"24",X"24",X"04",X"02",X"48",X"31",X"0A",X"FF",X"F2",
		X"4F",X"FF",X"42",X"42",X"42",X"42",X"03",X"07",X"0F",X"86",X"88",X"F8",X"B1",X"BB",X"8B",X"87",
		X"80",X"81",X"70",X"71",X"8B",X"87",X"80",X"F8",X"B1",X"BB",X"0F",X"86",X"88",X"03",X"07",X"0F",
		X"88",X"86",X"F8",X"1B",X"B0",X"8B",X"87",X"81",X"8B",X"70",X"70",X"81",X"87",X"80",X"F8",X"BB",
		X"10",X"0F",X"88",X"68",X"03",X"07",X"0F",X"88",X"68",X"F8",X"BB",X"1B",X"81",X"87",X"80",X"8B",
		X"70",X"70",X"8B",X"87",X"81",X"F8",X"1B",X"B0",X"0F",X"88",X"86",X"09",X"07",X"68",X"86",X"88",
		X"68",X"86",X"88",X"68",X"86",X"88",X"0B",X"B0",X"BB",X"0B",X"B0",X"BB",X"0B",X"B0",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"B0",X"BB",X"0B",X"B0",X"BB",
		X"0B",X"B0",X"BB",X"68",X"86",X"88",X"68",X"86",X"88",X"68",X"86",X"88",X"09",X"07",X"88",X"68",
		X"86",X"88",X"68",X"86",X"88",X"68",X"86",X"BB",X"0B",X"B0",X"BB",X"0B",X"B0",X"BB",X"0B",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"BB",X"0B",X"B0",X"BB",
		X"0B",X"B0",X"BB",X"0B",X"86",X"88",X"68",X"86",X"88",X"68",X"86",X"88",X"68",X"09",X"07",X"86",
		X"88",X"68",X"86",X"88",X"68",X"86",X"88",X"68",X"B0",X"BB",X"0B",X"B0",X"BB",X"0B",X"B0",X"BB",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"0B",X"B0",X"BB",
		X"0B",X"B0",X"BB",X"0B",X"B0",X"88",X"68",X"86",X"88",X"68",X"86",X"88",X"68",X"86",X"04",X"07",
		X"86",X"88",X"68",X"F0",X"B0",X"BB",X"1B",X"DF",X"00",X"08",X"78",X"B8",X"00",X"17",X"07",X"18",
		X"00",X"08",X"78",X"B8",X"B0",X"BB",X"1B",X"DF",X"86",X"88",X"68",X"F0",X"04",X"07",X"68",X"86",
		X"88",X"F0",X"0B",X"B1",X"BB",X"8F",X"00",X"08",X"78",X"18",X"00",X"07",X"07",X"B8",X"00",X"18",
		X"78",X"B8",X"BB",X"0B",X"B1",X"8F",X"88",X"68",X"88",X"F0",X"04",X"07",X"88",X"68",X"88",X"F0",
		X"BB",X"0B",X"B1",X"8F",X"00",X"18",X"78",X"B8",X"00",X"07",X"07",X"B8",X"00",X"08",X"78",X"18",
		X"0B",X"B1",X"BB",X"8F",X"68",X"86",X"88",X"F0",X"0C",X"06",X"00",X"00",X"0A",X"55",X"A0",X"AA",
		X"0A",X"55",X"A0",X"00",X"00",X"00",X"0A",X"55",X"A5",X"50",X"50",X"25",X"05",X"50",X"2A",X"AA",
		X"A0",X"00",X"02",X"20",X"02",X"25",X"A0",X"25",X"05",X"22",X"2A",X"55",X"55",X"00",X"00",X"25",
		X"02",X"50",X"00",X"25",X"0A",X"20",X"20",X"52",X"00",X"00",X"55",X"55",X"05",X"50",X"00",X"25",
		X"5A",X"50",X"50",X"55",X"00",X"00",X"AA",X"AA",X"0A",X"A0",X"00",X"55",X"5A",X"A0",X"A0",X"AA",
		X"00",X"00",X"0C",X"08",X"00",X"00",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BD",X"DD",X"DB",X"DD",X"DB",X"1D",X"BB",X"0B",X"00",X"BB",X"0B",X"D0",X"D1",X"11",X"1D",X"11",
		X"1B",X"1D",X"B1",X"B1",X"BB",X"D1",X"0B",X"10",X"00",X"D1",X"1D",X"10",X"1B",X"1D",X"01",X"B1",
		X"B1",X"10",X"0B",X"10",X"0D",X"1D",X"0D",X"DB",X"1B",X"1D",X"D1",X"B1",X"D1",X"00",X"0B",X"D0",
		X"DD",X"BB",X"BB",X"DD",X"DB",X"DB",X"DD",X"B1",X"BD",X"D0",X"00",X"00",X"DD",X"DD",X"DB",X"00",
		X"0B",X"D0",X"BD",X"BD",X"0B",X"DD",X"0B",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"D0",X"0C",X"08",X"0F",X"FF",X"F0",X"00",X"0F",X"66",X"F0",X"0F",X"F0",X"00",
		X"88",X"00",X"F6",X"66",X"68",X"00",X"06",X"DD",X"6F",X"06",X"DD",X"F8",X"66",X"F0",X"F1",X"60",
		X"F6",X"00",X"F1",X"0F",X"18",X"01",X"6D",X"66",X"61",X"F0",X"F1",X"6D",X"61",X"D0",X"B1",X"6D",
		X"1D",X"01",X"6F",X"6F",X"61",X"F0",X"F1",X"60",X"B6",X"10",X"D1",X"00",X"16",X"01",X"6B",X"FF",
		X"61",X"F0",X"F1",X"60",X"BD",X"10",X"DD",X"00",X"16",X"01",X"6B",X"0F",X"61",X"F0",X"FD",X"D1",
		X"1D",X"B0",X"BB",X"00",X"BB",X"06",X"60",X"00",X"66",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"F0",X"00",X"FF",X"00",X"0A",X"07",X"CC",X"4C",X"CC",X"44",X"4C",X"00",X"00",X"EE",
		X"04",X"C0",X"44",X"44",X"C9",X"4C",X"C9",X"40",X"00",X"4C",X"09",X"40",X"94",X"04",X"C9",X"C0",
		X"C9",X"4E",X"CE",X"4C",X"09",X"40",X"94",X"4C",X"C9",X"C0",X"C9",X"4C",X"4C",X"4C",X"04",X"C0",
		X"94",X"CC",X"09",X"4C",X"C4",X"94",X"94",X"4C",X"00",X"00",X"44",X"00",X"0C",X"44",X"CC",X"4E",
		X"04",X"CE",X"04",X"C0",X"CE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"40",X"08",X"07",
		X"88",X"88",X"00",X"99",X"00",X"04",X"40",X"00",X"80",X"00",X"09",X"00",X"90",X"40",X"04",X"00",
		X"88",X"80",X"09",X"00",X"90",X"40",X"04",X"00",X"00",X"08",X"09",X"00",X"90",X"40",X"04",X"00",
		X"00",X"08",X"09",X"00",X"90",X"40",X"04",X"00",X"80",X"08",X"09",X"00",X"90",X"40",X"04",X"00",
		X"08",X"80",X"00",X"99",X"00",X"04",X"40",X"00",X"0A",X"07",X"22",X"00",X"02",X"20",X"00",X"22",
		X"00",X"02",X"20",X"00",X"02",X"00",X"20",X"02",X"02",X"00",X"20",X"20",X"02",X"00",X"02",X"00",
		X"20",X"02",X"02",X"00",X"20",X"20",X"02",X"00",X"02",X"00",X"20",X"02",X"02",X"00",X"20",X"20",
		X"02",X"00",X"02",X"00",X"20",X"02",X"02",X"00",X"20",X"20",X"02",X"00",X"02",X"00",X"20",X"02",
		X"02",X"00",X"20",X"20",X"02",X"00",X"22",X"20",X"02",X"20",X"00",X"22",X"00",X"02",X"20",X"00",
		X"1E",X"B4",X"00",X"00",X"00",X"1F",X"6C",X"00",X"00",X"00",X"20",X"0C",X"00",X"00",X"00",X"20",
		X"C4",X"00",X"00",X"00",X"0A",X"0F",X"00",X"00",X"0C",X"71",X"37",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0C",X"C1",X"33",X"33",X"9C",X"00",X"00",X"00",X"00",X"00",X"CD",X"33",X"70",X"30",X"33",
		X"40",X"00",X"00",X"00",X"04",X"C3",X"73",X"43",X"23",X"43",X"C4",X"00",X"00",X"00",X"3E",X"CE",
		X"73",X"33",X"E3",X"9C",X"C7",X"4E",X"30",X"00",X"02",X"7C",X"C9",X"33",X"03",X"7C",X"EC",X"CA",
		X"97",X"30",X"00",X"0C",X"7C",X"73",X"97",X"CC",X"7E",X"C3",X"9C",X"70",X"00",X"0E",X"44",X"CE",
		X"EC",X"C4",X"7C",X"00",X"7E",X"00",X"00",X"00",X"C4",X"44",X"44",X"44",X"CE",X"00",X"00",X"00",
		X"00",X"00",X"8C",X"74",X"47",X"CC",X"E0",X"00",X"00",X"00",X"00",X"08",X"8F",X"F0",X"0F",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"08",X"FF",X"00",X"A8",X"F0",X"00",X"00",X"00",X"00",X"00",X"06",
		X"BF",X"00",X"0B",X"DB",X"00",X"00",X"00",X"00",X"00",X"BD",X"DE",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"1D",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"09",X"03",X"0B",
		X"02",X"0C",X"01",X"0D",X"00",X"10",X"01",X"12",X"03",X"12",X"03",X"11",X"04",X"0D",X"04",X"0C",
		X"03",X"0A",X"03",X"0A",X"03",X"0B",X"02",X"05",X"02",X"04",X"FF",X"FF",X"0A",X"0D",X"00",X"00",
		X"00",X"CD",X"13",X"97",X"E0",X"00",X"00",X"00",X"00",X"00",X"04",X"D3",X"33",X"33",X"BC",X"00",
		X"00",X"00",X"00",X"00",X"43",X"37",X"03",X"07",X"33",X"C0",X"00",X"00",X"00",X"04",X"C3",X"94",
		X"32",X"34",X"93",X"C4",X"00",X"00",X"00",X"44",X"CE",X"73",X"3C",X"33",X"7E",X"CC",X"40",X"00",
		X"03",X"EC",X"E4",X"C3",X"33",X"33",X"EC",X"EC",X"E3",X"00",X"37",X"90",X"C4",X"4C",X"93",X"9C",
		X"C7",X"C0",X"97",X"30",X"00",X"70",X"EC",X"44",X"CE",X"CC",X"4C",X"E0",X"70",X"00",X"00",X"00",
		X"08",X"E4",X"44",X"44",X"EF",X"00",X"00",X"00",X"00",X"00",X"0F",X"8E",X"C4",X"CE",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"00",X"08",X"80",X"00",X"00",X"00",X"00",X"00",X"0B",X"DB",
		X"F0",X"FB",X"DA",X"00",X"00",X"00",X"00",X"00",X"DD",X"DA",X"00",X"0A",X"DD",X"A0",X"00",X"00",
		X"06",X"0C",X"05",X"0D",X"04",X"0E",X"03",X"0F",X"02",X"10",X"01",X"11",X"00",X"12",X"02",X"10",
		X"05",X"0D",X"05",X"0D",X"06",X"0C",X"05",X"0D",X"04",X"0E",X"FF",X"FF",X"0A",X"0F",X"00",X"00",
		X"00",X"00",X"07",X"13",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"93",X"33",X"33",X"CE",
		X"00",X"00",X"00",X"00",X"00",X"C3",X"30",X"30",X"73",X"3D",X"C0",X"00",X"00",X"00",X"04",X"C3",
		X"43",X"23",X"43",X"93",X"CC",X"00",X"00",X"3E",X"47",X"CC",X"33",X"E3",X"33",X"7E",X"CE",X"90",
		X"37",X"9A",X"CC",X"EC",X"73",X"03",X"39",X"CC",X"79",X"00",X"7C",X"93",X"CE",X"74",X"C7",X"93",
		X"7C",X"CC",X"00",X"00",X"0E",X"70",X"0E",X"74",X"4C",X"EE",X"CC",X"4E",X"00",X"00",X"00",X"00",
		X"0E",X"C4",X"44",X"44",X"44",X"C0",X"00",X"00",X"00",X"00",X"00",X"EC",X"C7",X"44",X"7C",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"FF",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"A0",X"0F",X"F8",X"00",X"00",X"00",X"00",X"00",X"0B",X"DB",X"00",X"0F",X"B6",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"DD",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"ED",X"D0",X"00",X"09",X"0D",X"07",X"0F",X"06",X"10",X"05",X"11",X"02",X"12",X"00",X"11",
		X"00",X"0F",X"01",X"0F",X"05",X"0E",X"06",X"0E",X"08",X"0F",X"08",X"0F",X"07",X"0F",X"0D",X"10",
		X"0E",X"10",X"FF",X"FF",X"0B",X"0A",X"00",X"00",X"00",X"0C",X"D1",X"39",X"7E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"4D",X"33",X"33",X"3B",X"CC",X"00",X"00",X"00",X"03",X"E4",X"4C",X"33",
		X"39",X"39",X"33",X"3C",X"44",X"E3",X"00",X"37",X"9E",X"CE",X"39",X"43",X"23",X"49",X"3E",X"CE",
		X"77",X"30",X"99",X"73",X"E4",X"C7",X"33",X"E3",X"37",X"CC",X"E3",X"79",X"90",X"0C",X"70",X"C2",
		X"4C",X"33",X"03",X"3C",X"44",X"40",X"7C",X"00",X"00",X"00",X"C4",X"44",X"C9",X"39",X"C4",X"44",
		X"C0",X"00",X"00",X"00",X"00",X"0E",X"CC",X"4C",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AB",X"F8",X"88",X"FB",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"E0",X"00",X"ED",
		X"B0",X"00",X"00",X"00",X"07",X"0D",X"05",X"0F",X"01",X"13",X"00",X"14",X"00",X"14",X"01",X"13",
		X"04",X"10",X"05",X"0F",X"06",X"0E",X"06",X"0E",X"FF",X"FF",X"21",X"59",X"00",X"00",X"00",X"22",
		X"2E",X"00",X"00",X"00",X"22",X"E6",X"00",X"00",X"00",X"09",X"13",X"00",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"0A",X"B0",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"BB",X"BA",X"AA",X"00",X"00",X"00",X"00",X"00",X"C1",X"44",X"CC",X"CC",X"00",X"00",X"00",X"AB",
		X"BB",X"BB",X"BB",X"BA",X"AA",X"AA",X"A0",X"00",X"0A",X"D0",X"D0",X"00",X"00",X"00",X"EC",X"A0",
		X"00",X"00",X"E0",X"00",X"03",X"00",X"00",X"E0",X"00",X"00",X"00",X"AE",X"93",X"7E",X"79",X"9E",
		X"A0",X"00",X"00",X"0A",X"DA",X"73",X"33",X"33",X"7E",X"BB",X"00",X"00",X"0B",X"BA",X"AE",X"93",
		X"7E",X"11",X"EB",X"B0",X"00",X"0A",X"BB",X"AE",X"ED",X"11",X"19",X"11",X"BB",X"00",X"00",X"BB",
		X"BD",X"11",X"79",X"11",X"71",X"91",X"B0",X"00",X"0A",X"39",X"EC",X"CC",X"CC",X"CC",X"CE",X"30",
		X"00",X"00",X"B7",X"33",X"3A",X"AA",X"A0",X"33",X"70",X"00",X"00",X"AA",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"A0",X"0A",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"0A",
		X"D0",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"0A",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"0B",X"D0",X"00",X"00",X"09",X"09",X"06",X"0A",X"05",X"0B",X"04",X"0B",X"00",X"0E",
		X"01",X"0E",X"02",X"0C",X"02",X"0C",X"01",X"0D",X"01",X"0E",X"01",X"0F",X"02",X"10",X"03",X"10",
		X"04",X"10",X"04",X"06",X"05",X"0A",X"06",X"0A",X"05",X"0B",X"09",X"0C",X"FF",X"FF",X"08",X"12",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"0A",X"B0",X"00",X"00",
		X"00",X"00",X"0A",X"BB",X"BA",X"AA",X"00",X"00",X"00",X"00",X"C1",X"44",X"CC",X"CC",X"00",X"00",
		X"AB",X"BB",X"BB",X"BB",X"BA",X"AA",X"AA",X"A0",X"0A",X"D0",X"D0",X"00",X"00",X"00",X"EC",X"A0",
		X"00",X"E0",X"00",X"03",X"00",X"00",X"E0",X"00",X"00",X"BE",X"93",X"7E",X"73",X"9E",X"A0",X"00",
		X"0B",X"DA",X"73",X"33",X"33",X"7E",X"BA",X"00",X"AB",X"BA",X"AE",X"D1",X"1D",X"EA",X"AB",X"A0",
		X"BB",X"AA",X"D1",X"19",X"19",X"1D",X"AB",X"B0",X"0B",X"D1",X"97",X"11",X"17",X"91",X"1B",X"00",
		X"03",X"7C",X"C4",X"4C",X"CC",X"CE",X"73",X"00",X"00",X"73",X"33",X"AA",X"A3",X"33",X"70",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"A0",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"A0",X"AB",X"00",X"00",X"00",X"00",X"00",X"AB",X"A0",X"AB",X"A0",X"00",X"00",
		X"09",X"09",X"06",X"0A",X"05",X"0B",X"04",X"0B",X"00",X"0E",X"01",X"0E",X"02",X"0C",X"02",X"0C",
		X"01",X"0D",X"00",X"0E",X"00",X"0E",X"01",X"0D",X"01",X"0D",X"02",X"0C",X"12",X"00",X"05",X"09",
		X"05",X"09",X"04",X"0A",X"FF",X"FF",X"09",X"13",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AB",X"0A",X"B0",X"00",X"00",X"00",X"00",X"00",X"0A",X"BB",X"BA",
		X"AA",X"00",X"00",X"00",X"00",X"00",X"C1",X"44",X"CC",X"CC",X"00",X"00",X"00",X"AB",X"BB",X"BB",
		X"BB",X"BA",X"AA",X"AA",X"A0",X"00",X"0A",X"D0",X"D0",X"00",X"00",X"00",X"EC",X"A0",X"00",X"00",
		X"E0",X"00",X"03",X"00",X"00",X"E0",X"00",X"00",X"00",X"AE",X"93",X"7E",X"73",X"9E",X"A0",X"00",
		X"00",X"0B",X"AA",X"73",X"33",X"33",X"7E",X"AA",X"00",X"00",X"BA",X"E1",X"1E",X"93",X"7E",X"AA",
		X"BB",X"00",X"0B",X"B1",X"11",X"91",X"1D",X"EE",X"AA",X"BA",X"00",X"B1",X"19",X"71",X"11",X"79",
		X"1D",X"AB",X"B0",X"00",X"3E",X"CC",X"CC",X"CC",X"CC",X"E9",X"3A",X"00",X"00",X"73",X"30",X"AA",
		X"AA",X"33",X"97",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"DA",X"0A",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"BA",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"DB",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"0B",X"08",X"0C",X"07",X"0D",X"06",X"0D",X"02",X"10",X"03",X"10",X"04",
		X"0E",X"04",X"0E",X"03",X"0F",X"02",X"0F",X"01",X"0F",X"00",X"0E",X"00",X"0D",X"00",X"0C",X"0A",
		X"0C",X"06",X"0B",X"06",X"0A",X"05",X"0B",X"04",X"07",X"FF",X"FF",X"02",X"14",X"16",X"A2",X"04",
		X"10",X"10",X"51",X"02",X"00",X"10",X"9E",X"90",X"81",X"04",X"12",X"A2",X"08",X"60",X"41",X"0B",
		X"83",X"10",X"88",X"54",X"75",X"74",X"1E",X"83",X"94",X"42",X"B0",X"52",X"3C",X"0B",X"21",X"10",
		X"22",X"8E",X"0A",X"84",X"6B",X"A0",X"E0",X"12",X"96",X"92",X"A2",X"14",X"83",X"51",X"60",X"94",
		X"6D",X"2D",X"16",X"09",X"44",X"52",X"51",X"41",X"50",X"A5",X"64",X"1A",X"82",X"11",X"75",X"D4",
		X"42",X"80",X"C9",X"A9",X"29",X"81",X"08",X"52",X"92",X"9C",X"3A",X"3E",X"92",X"98",X"2A",X"16",
		X"AE",X"82",X"10",X"42",X"30",X"3A",X"10",X"AE",X"A2",X"12",X"82",X"11",X"34",X"E4",X"33",X"4F",
		X"42",X"74",X"E4",X"31",X"5D",X"0E",X"82",X"D1",X"21",X"D0",X"A5",X"65",X"10",X"88",X"12",X"8D",
		X"A5",X"21",X"EA",X"52",X"18",X"A5",X"21",X"BA",X"E8",X"60",X"08",X"26",X"0C",X"86",X"2A",X"A8",
		X"8F",X"82",X"50",X"3A",X"52",X"10",X"98",X"29",X"3D",X"31",X"0D",X"D5",X"51",X"1C",X"04",X"A0",
		X"65",X"A4",X"C3",X"E9",X"28",X"D0",X"52",X"32",X"92",X"87",X"6A",X"A8",X"8D",X"87",X"40",X"CF",
		X"4B",X"82",X"34",X"59",X"08",X"56",X"47",X"D2",X"21",X"95",X"54",X"46",X"43",X"A0",X"68",X"AD",
		X"14",X"BC",X"11",X"A2",X"28",X"22",X"A6",X"42",X"EA",X"A8",X"8B",X"87",X"40",X"9B",X"4A",X"82",
		X"D5",X"A2",X"12",X"A0",X"7D",X"4E",X"85",X"D4",X"51",X"15",X"0E",X"84",X"E9",X"30",X"EA",X"27",
		X"06",X"69",X"D0",X"4E",X"AC",X"42",X"6C",X"0E",X"AB",X"C6",X"24",X"42",X"AA",X"28",X"89",X"87",
		X"42",X"94",X"B8",X"55",X"1A",X"82",X"95",X"A3",X"12",X"60",X"85",X"58",X"84",X"42",X"06",X"F5",
		X"E2",X"92",X"A1",X"55",X"14",X"44",X"43",X"A3",X"E9",X"91",X"4B",X"47",X"A4",X"44",X"22",X"D0",
		X"BA",X"F1",X"6A",X"C4",X"26",X"C3",X"AA",X"C4",X"22",X"30",X"21",X"A5",X"43",X"AB",X"45",X"26",
		X"C2",X"6A",X"28",X"88",X"06",X"47",X"53",X"E2",X"97",X"8B",X"5E",X"21",X"19",X"84",X"D2",X"A2",
		X"51",X"38",X"65",X"58",X"84",X"4E",X"0E",X"53",X"A1",X"75",X"E2",X"13",X"E1",X"35",X"14",X"4E",
		X"0C",X"8E",X"AF",X"1C",X"9F",X"12",X"B4",X"52",X"37",X"1E",X"B4",X"62",X"91",X"28",X"A4",X"2A",
		X"AC",X"42",X"2B",X"05",X"28",X"AC",X"26",X"B4",X"52",X"21",X"09",X"A8",X"A2",X"68",X"54",X"75",
		X"78",X"C4",X"4A",X"25",X"58",X"A4",X"76",X"2D",X"68",X"84",X"88",X"94",X"56",X"13",X"56",X"64",
		X"3A",X"84",X"56",X"88",X"44",X"A1",X"35",X"14",X"4C",X"0A",X"8D",X"AF",X"14",X"8A",X"CE",X"AC",
		X"52",X"3F",X"12",X"AC",X"42",X"54",X"E8",X"BC",X"7A",X"1F",X"C6",X"AD",X"10",X"89",X"C2",X"6A",
		X"28",X"96",X"15",X"19",X"5E",X"29",X"17",X"9D",X"58",X"84",X"21",X"89",X"52",X"64",X"B8",X"94",
		X"5E",X"3D",X"0F",X"A3",X"55",X"88",X"45",X"21",X"35",X"14",X"4A",X"0A",X"8B",X"AF",X"14",X"8C",
		X"CE",X"AC",X"C8",X"45",X"12",X"9F",X"3A",X"33",X"1A",X"87",X"B1",X"6A",X"C4",X"22",X"90",X"AA",
		X"8A",X"24",X"85",X"45",X"D6",X"8A",X"46",X"A2",X"50",X"9E",X"74",X"F9",X"D6",X"8F",X"44",X"A2",
		X"D0",X"F2",X"25",X"58",X"84",X"56",X"13",X"55",X"44",X"80",X"A8",X"BA",X"D1",X"08",X"E4",X"E8",
		X"A4",X"52",X"4D",X"32",X"74",X"F9",X"D5",X"89",X"50",X"B5",X"11",X"8B",X"43",X"A8",X"95",X"62",
		X"11",X"68",X"4D",X"45",X"17",X"0A",X"8B",X"AD",X"10",X"8E",X"CE",X"89",X"46",X"25",X"D2",X"E7",
		X"4F",X"9D",X"58",X"95",X"4B",X"5C",X"88",X"45",X"A1",X"CC",X"EA",X"C4",X"22",X"D0",X"9A",X"AA",
		X"2C",X"15",X"17",X"5A",X"21",X"1D",X"89",X"44",X"63",X"13",X"69",X"53",X"A7",X"CE",X"AC",X"4A",
		X"A5",X"EE",X"44",X"22",X"D0",X"DE",X"25",X"59",X"91",X"78",X"4D",X"55",X"15",X"0A",X"8B",X"AD",
		X"10",X"8F",X"44",X"A2",X"11",X"C9",X"B4",X"A9",X"D3",X"E7",X"56",X"25",X"52",X"45",X"C8",X"84",
		X"5A",X"19",X"CC",X"F1",X"2A",X"CC",X"8B",X"C2",X"AA",X"28",X"A0",X"54",X"5D",X"68",X"84",X"7A",
		X"2D",X"10",X"8E",X"49",X"AA",X"7A",X"54",X"E9",X"F3",X"AB",X"0D",X"A8",X"44",X"22",X"D0",X"C6",
		X"67",X"89",X"56",X"64",X"62",X"13",X"55",X"45",X"02",X"22",X"EB",X"44",X"23",X"F1",X"69",X"F0",
		X"82",X"45",X"63",X"D2",X"A7",X"4F",X"9D",X"58",X"6D",X"52",X"21",X"16",X"85",X"D1",X"0A",X"4E",
		X"8E",X"42",X"AA",X"28",X"E1",X"51",X"55",X"A2",X"11",X"F8",X"D4",X"F8",X"49",X"7A",X"A7",X"A5",
		X"CE",X"9F",X"3A",X"D3",X"25",X"D5",X"22",X"31",X"68",X"59",X"10",X"A4",X"4A",X"37",X"0A",X"AA",
		X"A3",X"84",X"45",X"56",X"88",X"42",X"08",X"D4",X"F8",X"51",X"26",X"97",X"12",X"9F",X"3A",X"D1",
		X"09",X"35",X"CA",X"CC",X"9B",X"1A",X"85",X"11",X"4A",X"44",X"A3",X"70",X"BA",X"8A",X"38",X"44",
		X"55",X"58",X"84",X"20",X"84",X"53",X"A1",X"65",X"E9",X"93",X"A2",X"13",X"AF",X"10",X"BD",X"20",
		X"AC",X"C9",X"D1",X"E8",X"45",X"08",X"29",X"12",X"8D",X"C2",X"EA",X"A8",X"E1",X"11",X"35",X"62",
		X"11",X"28",X"B4",X"D8",X"55",X"36",X"1E",X"4D",X"9D",X"3E",X"74",X"88",X"79",X"58",X"84",X"E8",
		X"45",X"1E",X"8A",X"48",X"89",X"46",X"E1",X"95",X"14",X"70",X"88",X"9A",X"B1",X"08",X"84",X"22",
		X"97",X"0B",X"A7",X"43",X"09",X"D1",X"29",X"F3",X"A4",X"C3",X"8A",X"C4",X"27",X"C2",X"68",X"47",
		X"16",X"8D",X"C3",X"2A",X"A8",X"E1",X"11",X"35",X"62",X"13",X"E1",X"74",X"88",X"65",X"10",X"84",
		X"11",X"09",X"D1",X"09",X"D2",X"A1",X"A5",X"62",X"11",X"08",X"55",X"1D",X"84",X"51",X"B8",X"65",
		X"55",X"1C",X"22",X"26",X"AC",X"42",X"74",X"1B",X"A1",X"24",X"4A",X"7C",X"E9",X"90",X"B2",X"B1",
		X"08",X"94",X"2A",X"8D",X"42",X"A8",X"D4",X"36",X"AA",X"8E",X"11",X"13",X"56",X"21",X"3A",X"0D",
		X"D0",X"92",X"74",X"42",X"74",X"D8",X"51",X"59",X"91",X"48",X"4D",X"59",X"91",X"58",X"55",X"1A",
		X"86",X"D5",X"51",X"C2",X"22",X"6A",X"C4",X"27",X"C1",X"9A",X"12",X"44",X"A7",X"C4",X"A7",X"C7",
		X"2B",X"32",X"2D",X"08",X"AB",X"10",X"89",X"C2",X"A8",X"D4",X"36",X"AA",X"8E",X"11",X"13",X"56",
		X"21",X"08",X"21",X"14",X"23",X"89",X"44",X"27",X"42",X"E8",X"F5",X"62",X"11",X"28",X"55",X"1A",
		X"86",X"D5",X"51",X"C2",X"A2",X"6A",X"C4",X"21",X"0C",X"5A",X"3D",X"32",X"D1",X"28",X"8C",X"E8",
		X"5F",X"1A",X"AC",X"42",X"25",X"0A",X"A3",X"10",X"EA",X"AA",X"38",X"54",X"4D",X"68",X"84",X"20",
		X"8B",X"47",X"22",X"16",X"89",X"44",X"62",X"50",X"BE",X"35",X"59",X"91",X"28",X"55",X"17",X"87",
		X"D5",X"51",X"40",X"A8",X"9A",X"D1",X"08",X"41",X"3A",X"37",X"14",X"B4",X"4A",X"25",X"12",X"86",
		X"11",X"6A",X"CC",X"89",X"42",X"A8",X"A4",X"11",X"AA",X"A2",X"A1",X"11",X"55",X"A3",X"91",X"C9",
		X"D1",X"A8",X"A5",X"62",X"D1",X"28",X"B4",X"31",X"89",X"56",X"64",X"4A",X"13",X"44",X"60",X"A5",
		X"55",X"16",X"08",X"8A",X"AF",X"14",X"8E",X"4E",X"8C",X"45",X"2D",X"12",X"8A",X"45",X"A1",X"94",
		X"4A",X"29",X"09",X"A7",X"C1",X"6A",X"AA",X"2C",X"15",X"15",X"44",X"A3",X"13",X"E7",X"47",X"A2",
		X"51",X"48",X"D4",X"33",X"89",X"44",X"E1",X"34",X"E8",X"2D",X"55",X"45",X"82",X"A3",X"28",X"9C",
		X"42",X"74",X"E8",X"E4",X"5A",X"2B",X"1A",X"8E",X"CC",X"8C",X"44",X"A2",X"50",X"8A",X"74",X"16",
		X"AA",X"A2",X"C1",X"50",X"85",X"10",X"88",X"4D",X"9D",X"1A",X"8B",X"45",X"A3",X"D1",X"E8",X"84",
		X"5E",X"74",X"46",X"13",X"4D",X"82",X"D5",X"54",X"54",X"2A",X"1C",X"AD",X"32",X"6C",X"E8",X"BC",
		X"7A",X"2D",X"0C",X"A2",X"91",X"AA",X"C4",X"22",X"D1",X"28",X"84",X"26",X"99",X"05",X"AA",X"A8",
		X"A0",X"54",X"3D",X"56",X"64",X"D9",X"D1",X"68",X"F4",X"20",X"8B",X"44",X"A3",X"D5",X"88",X"45",
		X"A7",X"4F",X"84",X"D3",X"60",X"AD",X"55",X"14",X"08",X"8F",X"A4",X"43",X"2A",X"CC",X"9B",X"3A",
		X"2B",X"08",X"A1",X"14",X"4A",X"23",X"08",X"AB",X"10",X"8A",X"CE",X"9F",X"09",X"A6",X"41",X"5A",
		X"AA",X"38",X"54",X"6D",X"32",X"15",X"56",X"64",X"D9",X"D1",X"58",X"F4",X"24",X"89",X"44",X"21",
		X"35",X"62",X"11",X"49",X"D3",X"A1",X"34",X"C8",X"2B",X"55",X"47",X"0A",X"8C",X"AD",X"1C",X"AC",
		X"22",X"AC",X"C9",X"D3",X"A2",X"90",X"8A",X"12",X"44",X"A2",X"30",X"9A",X"B1",X"08",X"9C",X"E9",
		X"D0",X"9A",X"5C",X"32",X"A2",X"22",X"B2",X"8A",X"A3",X"2B",X"46",X"24",X"46",X"AB",X"32",X"7C",
		X"E8",X"A4",X"7A",X"13",X"44",X"A2",X"10",X"AA",X"B1",X"08",X"94",X"E9",X"B0",X"AA",X"5C",X"2E",
		X"9A",X"A2",X"A8",X"BA",X"D1",X"09",X"91",X"28",X"A4",X"E8",X"9C",X"22",X"84",X"F3",X"A2",X"10",
		X"BA",X"B1",X"08",X"8C",X"E9",X"B0",X"AA",X"54",X"2E",X"98",X"A2",X"88",X"CA",X"B1",X"08",X"41",
		X"12",X"89",X"C7",X"A1",X"44",X"E8",X"84",X"32",X"AC",X"42",X"21",X"3A",X"64",X"2E",X"93",X"0B",
		X"AA",X"A2",X"88",X"BA",X"B1",X"08",X"43",X"3A",X"D3",X"27",X"C7",X"A1",X"44",X"E8",X"84",X"36",
		X"AC",X"42",X"7C",X"E9",X"70",X"DA",X"F0",X"BA",X"AA",X"28",X"8B",X"AB",X"10",X"84",X"11",X"2A",
		X"CC",X"9F",X"1E",X"85",X"33",X"A2",X"10",X"EA",X"B1",X"09",X"B1",X"29",X"70",X"EA",X"B0",X"BA",
		X"AA",X"28",X"8B",X"AB",X"32",X"10",X"C4",X"AB",X"32",X"74",X"22",X"85",X"11",X"28",X"84",X"3E",
		X"AC",X"42",X"F1",X"0A",X"44",X"A5",X"C1",X"AA",X"AA",X"28",X"8B",X"AB",X"32",X"10",X"45",X"AB",
		X"32",X"74",X"7A",X"12",X"CC",X"A4",X"4A",X"21",X"04",X"6A",X"C2",X"4A",X"44",X"A6",X"41",X"9A",
		X"AA",X"28",X"8B",X"AB",X"32",X"39",X"32",X"91",X"AA",X"CC",X"9B",X"08",X"A1",X"24",X"42",X"93",
		X"A6",X"CC",X"AC",X"12",X"A6",X"44",X"A6",X"47",X"A4",X"43",X"AA",X"A8",X"AA",X"2A",X"AC",X"C8",
		X"D4",X"42",X"B1",X"AA",X"C4",X"25",X"C2",X"28",X"45",X"18",X"A4",X"4A",X"64",X"CA",X"C1",X"5A",
		X"4C",X"4A",X"6C",X"6A",X"5C",X"32",X"AA",X"8A",X"A2",X"AB",X"4C",X"8C",X"44",X"2B",X"1E",X"AC",
		X"42",X"5C",X"22",X"8A",X"41",X"32",X"91",X"2B",X"4C",X"B4",X"42",X"B0",X"7A",X"9B",X"1A",X"AC",
		X"62",X"F0",X"AA",X"AA",X"38",X"54",X"55",X"1A",X"8A",X"56",X"11",X"56",X"21",X"2A",X"11",X"44",
		X"E1",X"24",X"F8",X"D5",X"E3",X"15",X"83",X"74",X"46",X"2D",X"58",X"A4",X"A8",X"55",X"55",X"1C",
		X"2A",X"2A",X"BC",X"C8",X"94",X"52",X"D0",X"9A",X"D1",X"09",X"30",X"8A",X"25",X"14",X"89",X"42",
		X"69",X"90",X"72",X"88",X"45",X"AB",X"14",X"97",X"0B",X"A8",X"A2",X"81",X"51",X"54",X"5A",X"29",
		X"68",X"5D",X"68",X"87",X"99",X"58",X"4D",X"10",X"8A",X"4A",X"82",X"B4",X"98",X"3D",X"4E",X"8D",
		X"52",X"29",X"36",X"15",X"55",X"45",X"02",X"A2",X"E8",X"94",X"62",X"D0",X"DA",X"6C",X"2A",X"9B",
		X"14",X"B4",X"1C",X"AD",X"0F",X"AC",X"84",X"29",X"71",X"EA",X"45",X"27",X"42",X"AA",X"A8",X"A8",
		X"54",X"5D",X"18",X"87",X"D2",X"E1",X"75",X"E6",X"56",X"29",X"68",X"17",X"52",X"50",X"85",X"78",
		X"4D",X"48",X"84",X"F8",X"55",X"55",X"15",X"0C",X"8B",X"A2",X"90",X"4E",X"93",X"0D",X"A4",X"45",
		X"2D",X"02",X"FA",X"5A",X"1B",X"A9",X"10",X"9F",X"0A",X"AA",X"A2",X"C1",X"51",X"B4",X"C8",X"37",
		X"56",X"08",X"53",X"20",X"61",X"59",X"30",X"54",X"35",X"52",X"21",X"3E",X"15",X"55",X"45",X"C2",
		X"A3",X"69",X"50",X"2F",X"A4",X"40",X"CA",X"AA",X"20",X"2A",X"19",X"A9",X"10",X"9F",X"0A",X"AA",
		X"A2",X"40",X"54",X"75",X"68",X"0C",X"D5",X"51",X"41",X"90",X"BD",X"58",X"84",X"D8",X"5D",X"55",
		X"12",X"42",X"A0",X"50",X"A2",X"C8",X"4A",X"AA",X"30",X"32",X"17",X"AB",X"10",X"99",X"0B",X"A8",
		X"A2",X"50",X"54",X"3B",X"59",X"05",X"94",X"75",X"1D",X"55",X"1E",X"19",X"0B",X"53",X"E1",X"75",
		X"54",X"4B",X"0C",X"86",X"69",X"68",X"28",X"A4",X"21",X"10",X"5A",X"2A",X"B2",X"11",X"0E",X"85",
		X"69",X"B0",X"CA",X"8A",X"26",X"06",X"42",X"F4",X"D4",X"25",X"59",X"09",X"56",X"43",X"00",X"94",
		X"D5",X"D0",X"A0",X"74",X"2B",X"4A",X"86",X"55",X"51",X"34",X"3A",X"10",X"A5",X"27",X"0E",X"8F",
		X"A4",X"23",X"69",X"08",X"74",X"1C",X"85",X"C1",X"68",X"46",X"B4",X"36",X"AA",X"89",X"C0",X"84",
		X"6D",X"25",X"16",X"08",X"45",X"D2",X"D1",X"54",X"84",X"10",X"02",X"90",X"E0",X"31",X"0D",X"D5",
		X"51",X"10",X"04",X"22",X"29",X"48",X"F0",X"22",X"98",X"10",X"96",X"BA",X"04",X"A0",X"4A",X"18",
		X"AA",X"A2",X"24",X"04",X"10",X"B0",X"35",X"12",X"0C",X"40",X"9E",X"1D",X"0B",X"55",X"51",X"14",
		X"05",X"A1",X"B0",X"4A",X"30",X"14",X"81",X"48",X"32",X"14",X"AA",X"A2",X"09",X"21",X"90",X"2A",
		X"86",X"42",X"55",X"54",X"40",X"A2",X"0C",X"8E",X"AC",X"A2",X"05",X"18",X"74",X"55",X"75",X"10",
		X"29",X"00",X"8A",X"88",X"14",X"C0",X"D5",X"18",X"00",X"2B",X"0D",X"00",X"00",X"00",X"2B",X"9F",
		X"00",X"00",X"00",X"2C",X"0D",X"00",X"00",X"00",X"2C",X"63",X"00",X"00",X"00",X"0C",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"12",
		X"70",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"92",X"99",X"E0",X"07",X"9E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"2E",X"72",X"97",X"E0",X"00",X"E7",X"97",X"00",X"79",
		X"77",X"92",X"7E",X"92",X"7E",X"79",X"99",X"99",X"97",X"00",X"90",X"00",X"00",X"00",X"00",X"E9",
		X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"29",X"99",X"7E",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",
		X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"12",X"27",
		X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"92",X"22",X"90",X"00",X"09",X"00",X"00",X"00",X"00",
		X"72",X"E7",X"92",X"E7",X"90",X"00",X"00",X"00",X"00",X"07",X"92",X"E9",X"99",X"E0",X"00",X"90",
		X"90",X"79",X"77",X"77",X"2E",X"77",X"99",X"97",X"00",X"79",X"7E",X"00",X"07",X"79",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"0E",X"97",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"79",X"70",X"00",X"00",X"00",X"00",X"07",X"0C",X"72",
		X"7E",X"00",X"00",X"00",X"00",X"00",X"02",X"12",X"70",X"00",X"00",X"00",X"00",X"E9",X"2E",X"27",
		X"00",X"00",X"00",X"00",X"07",X"99",X"E2",X"70",X"00",X"00",X"00",X"00",X"79",X"2E",X"27",X"00",
		X"00",X"00",X"00",X"07",X"99",X"72",X"09",X"00",X"00",X"00",X"0E",X"72",X"E7",X"90",X"00",X"00",
		X"00",X"07",X"09",X"70",X"99",X"00",X"20",X"90",X"07",X"02",X"70",X"07",X"99",X"E0",X"07",X"9E",
		X"09",X"70",X"00",X"00",X"00",X"00",X"00",X"09",X"E0",X"00",X"00",X"00",X"00",X"00",X"27",X"00",
		X"00",X"00",X"00",X"09",X"04",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"29",X"7E",X"00",X"00",X"00",X"00",X"00",X"E7",X"97",X"EE",X"79",X"97",X"99",X"99",X"77",X"70",
		X"00",X"00",X"09",X"0E",X"E7",X"7E",X"00",X"00",X"00",X"04",X"05",X"00",X"D1",X"00",X"00",X"00",
		X"11",X"D0",X"00",X"10",X"17",X"91",X"B0",X"11",X"19",X"91",X"10",X"01",X"10",X"01",X"00",X"02",
		X"03",X"02",X"04",X"00",X"06",X"00",X"06",X"01",X"05",X"FF",X"FF",X"2C",X"FB",X"01",X"80",X"FC",
		X"2C",X"FB",X"FE",X"00",X"FA",X"2C",X"FB",X"FA",X"80",X"F6",X"2C",X"FB",X"F7",X"00",X"FA",X"2C",
		X"FB",X"F4",X"80",X"FD",X"2C",X"FB",X"F7",X"00",X"01",X"2C",X"FB",X"FA",X"80",X"04",X"2C",X"FB",
		X"FE",X"00",X"01",X"2C",X"FB",X"FD",X"00",X"FC",X"2C",X"FB",X"00",X"80",X"FA",X"2C",X"FB",X"04",
		X"00",X"F6",X"2C",X"FB",X"07",X"80",X"FA",X"2C",X"FB",X"0C",X"00",X"FD",X"2C",X"FB",X"07",X"80",
		X"01",X"2C",X"FB",X"04",X"00",X"05",X"2C",X"FB",X"00",X"80",X"01",X"08",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"79",X"00",X"00",X"09",X"79",X"00",X"00",X"07",X"00",X"70",
		X"00",X"00",X"70",X"00",X"00",X"09",X"00",X"7E",X"99",X"77",X"77",X"70",X"00",X"07",X"EE",X"7E",
		X"EE",X"EE",X"EE",X"E0",X"00",X"00",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"0B",X"01",X"0A",X"01",X"0C",X"01",X"0C",X"02",X"03",X"FF",X"FF",X"04",X"26",X"00",X"00",X"DD",
		X"00",X"00",X"0D",X"D8",X"00",X"00",X"DD",X"88",X"00",X"0D",X"D8",X"88",X"00",X"DD",X"88",X"A8",
		X"00",X"D8",X"8F",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",
		X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",
		X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"A8",
		X"00",X"D8",X"AA",X"88",X"00",X"D8",X"A8",X"88",X"00",X"D8",X"89",X"A8",X"00",X"D8",X"99",X"F8",
		X"00",X"D8",X"A7",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",
		X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"F8",
		X"00",X"D8",X"AF",X"F8",X"00",X"D8",X"AF",X"A8",X"00",X"D8",X"AA",X"88",X"00",X"D8",X"A8",X"8B",
		X"00",X"D8",X"88",X"B0",X"00",X"D8",X"8B",X"00",X"00",X"D8",X"B0",X"00",X"00",X"DB",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"09",X"26",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0D",X"DB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"EE",X"F8",X"88",X"88",X"88",
		X"88",X"00",X"0D",X"DE",X"EE",X"F8",X"88",X"88",X"88",X"88",X"00",X"DD",X"EE",X"EE",X"F8",X"AF",
		X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",
		X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",
		X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",
		X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",
		X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",
		X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",
		X"EE",X"F8",X"AA",X"AA",X"AA",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"88",X"88",X"88",X"88",X"00",
		X"DE",X"EE",X"EE",X"F8",X"88",X"88",X"89",X"98",X"00",X"DE",X"EE",X"EE",X"F8",X"88",X"88",X"8F",
		X"A8",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",
		X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DC",X"EE",X"EE",
		X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DC",
		X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"CE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",
		X"00",X"DC",X"EE",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"CE",X"EE",X"F8",X"AF",X"FF",
		X"FF",X"88",X"00",X"DC",X"EC",X"EE",X"F8",X"AF",X"FF",X"FF",X"88",X"00",X"DE",X"CE",X"EE",X"F8",
		X"AA",X"AA",X"AA",X"88",X"00",X"DC",X"EC",X"EE",X"F8",X"88",X"88",X"88",X"88",X"00",X"DE",X"CE",
		X"CE",X"F8",X"88",X"88",X"88",X"88",X"00",X"DC",X"EC",X"CB",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DC",X"CE",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"DC",X"EB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DC",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"26",X"DD",
		X"00",X"00",X"00",X"8D",X"D0",X"00",X"00",X"88",X"DD",X"00",X"00",X"88",X"8D",X"D0",X"00",X"8A",
		X"88",X"DD",X"00",X"8A",X"F8",X"8D",X"00",X"8A",X"FA",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",
		X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",
		X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",
		X"FF",X"8D",X"00",X"88",X"AF",X"8D",X"00",X"88",X"8A",X"8D",X"00",X"8A",X"98",X"8D",X"00",X"8A",
		X"99",X"8D",X"00",X"8A",X"7A",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",
		X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",
		X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"8A",X"FF",X"8D",X"00",X"88",X"AF",X"8D",X"00",X"B8",
		X"8A",X"8D",X"00",X"0B",X"88",X"8D",X"00",X"00",X"B8",X"8D",X"00",X"00",X"0B",X"8D",X"00",X"00",
		X"00",X"BD",X"00",X"00",X"00",X"0B",X"00",X"09",X"26",X"00",X"00",X"00",X"00",X"00",X"DD",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"D0",X"00",X"00",X"88",X"88",X"88",X"88",X"8F",
		X"EE",X"DD",X"00",X"00",X"88",X"88",X"88",X"88",X"8F",X"EE",X"ED",X"D0",X"00",X"88",X"AF",X"FF",
		X"FF",X"8F",X"EE",X"EE",X"DD",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",
		X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",
		X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",
		X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",
		X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",
		X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",
		X"88",X"AA",X"AA",X"AA",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"88",X"88",X"88",X"8F",X"EE",X"EE",
		X"ED",X"00",X"89",X"98",X"88",X"88",X"8F",X"EE",X"EE",X"ED",X"00",X"8A",X"F8",X"88",X"88",X"8F",
		X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",
		X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",X"00",X"88",
		X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"CD",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"ED",
		X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"CD",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",
		X"EC",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"EE",X"CD",X"00",X"88",X"AF",X"FF",X"FF",
		X"8F",X"EE",X"EC",X"ED",X"00",X"88",X"AF",X"FF",X"FF",X"8F",X"EE",X"CE",X"CD",X"00",X"88",X"AA",
		X"AA",X"AA",X"8F",X"EE",X"EC",X"ED",X"00",X"88",X"88",X"88",X"88",X"8F",X"EE",X"CE",X"CD",X"00",
		X"88",X"88",X"88",X"88",X"8F",X"EC",X"EC",X"ED",X"00",X"00",X"00",X"00",X"00",X"00",X"BC",X"CE",
		X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"EC",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BE",X"CD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"CD",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"10",
		X"03",X"00",X"00",X"00",X"FD",X"DD",X"DF",X"FF",X"FF",X"FF",X"FF",X"DD",X"DD",X"DF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FD",X"D8",X"88",X"88",X"88",X"88",X"8D",X"DF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"1D",X"1D",X"1D",X"D0",X"0D",X"D1",X"D1",X"D1",X"00",X"00",X"00",
		X"00",X"10",X"07",X"00",X"00",X"00",X"FD",X"DD",X"DF",X"FF",X"FF",X"FF",X"FF",X"FD",X"DD",X"DF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"FD",X"D8",X"88",X"88",X"88",X"88",X"8D",X"DF",X"81",
		X"00",X"00",X"00",X"00",X"00",X"00",X"1D",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"D1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"10",X"05",X"00",X"00",X"01",X"FD",X"DD",X"DF",X"FF",X"FF",X"FF",X"FF",X"FD",
		X"DD",X"DF",X"10",X"00",X"00",X"00",X"00",X"1D",X"D8",X"FD",X"D8",X"88",X"88",X"88",X"88",X"8D",
		X"DF",X"8D",X"D1",X"00",X"00",X"00",X"01",X"DD",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"DD",X"10",X"00",X"00",X"1D",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"D1",X"00",X"01",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"10",X"32",X"2E",X"05",X"00",X"07",X"32",X"5A",X"05",X"00",X"06",X"32",
		X"94",X"04",X"00",X"05",X"32",X"DE",X"01",X"F4",X"01",X"33",X"7C",X"00",X"00",X"04",X"06",X"05",
		X"00",X"05",X"E5",X"00",X"00",X"00",X"00",X"E5",X"94",X"19",X"00",X"00",X"00",X"44",X"44",X"1E",
		X"90",X"00",X"0D",X"81",X"4E",X"E9",X"91",X"E0",X"91",X"D8",X"EE",X"97",X"E7",X"90",X"03",X"05",
		X"02",X"07",X"02",X"08",X"01",X"0A",X"00",X"0A",X"FF",X"FF",X"07",X"06",X"00",X"07",X"9E",X"DE",
		X"00",X"00",X"00",X"00",X"09",X"5E",X"54",X"90",X"00",X"00",X"00",X"9E",X"59",X"D4",X"89",X"E0",
		X"00",X"09",X"C4",X"44",X"DA",X"E8",X"40",X"00",X"EC",X"D8",X"14",X"EE",X"99",X"E9",X"E0",X"C9",
		X"1D",X"8E",X"E9",X"9E",X"79",X"C0",X"03",X"07",X"03",X"08",X"02",X"0A",X"01",X"0A",X"00",X"0C",
		X"00",X"0C",X"FF",X"FF",X"08",X"07",X"00",X"00",X"0E",X"9A",X"D0",X"00",X"00",X"00",X"00",X"00",
		X"09",X"ED",X"9C",X"E0",X"00",X"00",X"00",X"00",X"95",X"E5",X"49",X"6E",X"00",X"00",X"00",X"79",
		X"E5",X"9D",X"4E",X"E6",X"E0",X"00",X"00",X"9E",X"C4",X"4D",X"AE",X"6E",X"6C",X"00",X"01",X"CE",
		X"81",X"4E",X"E9",X"9E",X"9E",X"00",X"1E",X"91",X"D8",X"EE",X"99",X"EE",X"91",X"00",X"05",X"08",
		X"05",X"0A",X"04",X"0B",X"02",X"0C",X"02",X"0D",X"01",X"0D",X"00",X"0D",X"FF",X"FF",X"0C",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"04",X"C0",X"00",X"00",X"00",X"0D",
		X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"90",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"00",X"00",X"00",X"99",X"E0",X"00",X"02",X"70",X"0E",X"29",X"50",X"00",X"0F",
		X"60",X"09",X"00",X"00",X"00",X"00",X"20",X"07",X"9E",X"5C",X"0C",X"E9",X"69",X"E0",X"00",X"00",
		X"90",X"00",X"00",X"C9",X"C4",X"44",X"DA",X"E6",X"E6",X"90",X"00",X"00",X"00",X"00",X"00",X"DC",
		X"E8",X"14",X"EE",X"99",X"E9",X"EC",X"00",X"60",X"00",X"00",X"0D",X"E9",X"1D",X"8E",X"E9",X"9E",
		X"E9",X"C1",X"00",X"00",X"0D",X"0D",X"08",X"10",X"05",X"10",X"06",X"07",X"15",X"16",X"09",X"16",
		X"03",X"13",X"04",X"12",X"00",X"12",X"06",X"16",X"05",X"13",X"FF",X"FF",X"0F",X"08",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"BD",X"DB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E0",X"00",X"0E",X"9A",X"D0",X"00",X"00",X"00",X"A1",X"00",X"00",X"00",X"50",X"00",X"EE",
		X"00",X"00",X"09",X"EC",X"9C",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E7",X"E0",X"00",
		X"00",X"95",X"E5",X"49",X"8E",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"4C",X"00",X"00",X"79",
		X"E5",X"9D",X"4E",X"E6",X"E0",X"00",X"EC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"C4",
		X"4D",X"AE",X"6E",X"6C",X"00",X"0E",X"7E",X"00",X"00",X"00",X"7E",X"00",X"01",X"CE",X"81",X"4E",
		X"E9",X"9E",X"9E",X"00",X"00",X"E7",X"90",X"90",X"09",X"70",X"00",X"1E",X"21",X"D8",X"EE",X"99",
		X"EE",X"91",X"00",X"00",X"0E",X"20",X"1C",X"1C",X"20",X"00",X"20",X"00",X"15",X"19",X"08",X"19",
		X"02",X"12",X"04",X"1C",X"04",X"19",X"0A",X"1B",X"04",X"1C",X"00",X"1C",X"FF",X"FF",X"34",X"1D",
		X"00",X"00",X"00",X"35",X"01",X"00",X"00",X"02",X"35",X"D7",X"00",X"00",X"FE",X"0C",X"10",X"00",
		X"00",X"00",X"0B",X"AD",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"DB",
		X"BB",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BD",X"BD",X"BB",X"AB",X"BA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EB",X"BB",X"BB",X"BB",X"BB",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"DB",X"BA",X"BA",X"AA",X"BA",X"00",X"00",X"00",X"00",X"0A",X"BA",X"EA",X"BB",
		X"AA",X"AA",X"DD",X"AB",X"AA",X"00",X"00",X"00",X"AD",X"BA",X"BA",X"BB",X"AD",X"1D",X"11",X"1A",
		X"AB",X"A0",X"00",X"00",X"DB",X"BB",X"BB",X"AB",X"A1",X"11",X"DB",X"CD",X"BA",X"BA",X"00",X"00",
		X"AB",X"BB",X"BB",X"BB",X"AD",X"1C",X"AB",X"0D",X"AA",X"AA",X"00",X"00",X"EA",X"DB",X"BB",X"BB",
		X"AA",X"D0",X"AA",X"BA",X"AB",X"AB",X"00",X"0A",X"BA",X"BB",X"BB",X"BB",X"BB",X"AA",X"BB",X"BA",
		X"BA",X"AA",X"00",X"AB",X"AB",X"BB",X"AB",X"BB",X"BB",X"BB",X"BA",X"AB",X"AB",X"AE",X"00",X"DA",
		X"BB",X"BA",X"BA",X"BA",X"BB",X"BB",X"AB",X"AA",X"AA",X"A0",X"00",X"EA",X"BA",X"BA",X"EA",X"EB",
		X"AB",X"AB",X"AA",X"AA",X"AE",X"00",X"00",X"0E",X"AA",X"AE",X"00",X"EA",X"AA",X"BA",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"07",
		X"0B",X"06",X"0D",X"06",X"0F",X"06",X"10",X"07",X"11",X"03",X"13",X"02",X"14",X"02",X"15",X"02",
		X"15",X"02",X"15",X"01",X"15",X"00",X"15",X"00",X"14",X"00",X"13",X"01",X"0E",X"09",X"0D",X"FF",
		X"FF",X"0D",X"0E",X"00",X"00",X"00",X"00",X"00",X"AD",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"BB",X"BB",X"AD",X"BE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"ED",X"BB",X"AB",X"AA",X"AB",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"BB",X"BA",
		X"AA",X"AD",X"DB",X"AA",X"00",X"00",X"00",X"00",X"00",X"ED",X"AA",X"DB",X"BA",X"D1",X"DB",X"11",
		X"AA",X"00",X"00",X"00",X"00",X"0E",X"DB",X"DB",X"BB",X"AA",X"11",X"1B",X"11",X"DA",X"A0",X"00",
		X"00",X"00",X"0A",X"BD",X"BB",X"BB",X"BA",X"D1",X"1A",X"BD",X"DA",X"AA",X"00",X"00",X"00",X"0E",
		X"AB",X"BB",X"BA",X"BA",X"AD",X"DA",X"AB",X"AA",X"BA",X"A0",X"00",X"0A",X"DB",X"DB",X"BB",X"BB",
		X"BB",X"BA",X"AB",X"BA",X"BB",X"AA",X"AE",X"00",X"AB",X"BB",X"BB",X"BA",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"AB",X"AA",X"AA",X"00",X"DB",X"DB",X"BB",X"AA",X"AD",X"BB",X"BB",X"BA",X"AA",X"BA",X"BA",
		X"AA",X"00",X"EA",X"BA",X"BB",X"EA",X"EA",X"BB",X"BA",X"BA",X"AE",X"AA",X"AB",X"AE",X"00",X"0E",
		X"AA",X"AE",X"00",X"0E",X"AA",X"BB",X"AA",X"E0",X"EA",X"AA",X"E0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"AA",X"AE",X"00",X"00",X"00",X"00",X"00",X"0A",X"0D",X"09",X"11",X"08",X"12",X"07",
		X"13",X"04",X"13",X"03",X"14",X"03",X"15",X"03",X"16",X"01",X"17",X"00",X"17",X"00",X"17",X"00",
		X"17",X"01",X"16",X"0B",X"0F",X"FF",X"FF",X"0B",X"10",X"00",X"00",X"00",X"0A",X"BB",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"DB",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"DB",X"BD",X"BA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"BB",
		X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"AB",X"BA",X"BA",X"AA",X"AB",X"A0",X"00",X"00",
		X"00",X"0A",X"BE",X"AD",X"BA",X"AA",X"DD",X"AB",X"AB",X"00",X"00",X"00",X"DB",X"DA",X"BB",X"AD",
		X"DB",X"0C",X"1A",X"AA",X"A0",X"00",X"0E",X"BB",X"BD",X"BB",X"A1",X"C0",X"B1",X"11",X"BB",X"A0",
		X"00",X"0A",X"AD",X"BB",X"BB",X"AD",X"11",X"AB",X"DD",X"AA",X"E0",X"00",X"0E",X"BB",X"BB",X"BB",
		X"AA",X"1D",X"AA",X"BA",X"BA",X"BA",X"00",X"AB",X"AB",X"BB",X"BB",X"BB",X"AA",X"BB",X"AB",X"AA",
		X"AB",X"00",X"BA",X"BB",X"BB",X"BA",X"BB",X"BB",X"BB",X"AA",X"AB",X"AA",X"00",X"EB",X"AB",X"DB",
		X"BB",X"BB",X"BB",X"BA",X"BA",X"BA",X"AE",X"00",X"0A",X"AA",X"BA",X"BA",X"BA",X"BA",X"BA",X"AA",
		X"AA",X"A0",X"00",X"00",X"EA",X"AA",X"EE",X"EB",X"AB",X"AB",X"EA",X"AE",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EA",X"AA",X"AE",X"00",X"00",X"00",X"00",X"07",X"0A",X"06",X"0B",X"06",X"0C",X"06",
		X"0E",X"06",X"10",X"03",X"11",X"02",X"12",X"01",X"12",X"01",X"12",X"01",X"13",X"00",X"13",X"00",
		X"13",X"00",X"13",X"01",X"12",X"02",X"11",X"08",X"0D",X"FF",X"FF",X"90",X"24",X"14",X"20",X"01",
		X"90",X"24",X"14",X"20",X"01",X"80",X"24",X"40",X"01",X"90",X"24",X"30",X"01",X"20",X"14",X"60",
		X"44",X"10",X"01",X"20",X"24",X"40",X"54",X"10",X"01",X"20",X"24",X"40",X"54",X"10",X"01",X"20",
		X"44",X"20",X"54",X"10",X"01",X"74",X"64",X"10",X"01",X"10",X"A4",X"30",X"01",X"10",X"A4",X"30",
		X"01",X"10",X"A4",X"30",X"01",X"40",X"6C",X"40",X"00",X"10",X"5C",X"01",X"6C",X"01",X"3C",X"14",
		X"3C",X"01",X"2C",X"34",X"2C",X"01",X"2C",X"34",X"2C",X"01",X"3C",X"14",X"3C",X"01",X"10",X"5C",
		X"01",X"10",X"3C",X"00",X"E0",X"01",X"E0",X"01",X"E0",X"01",X"E0",X"01",X"A0",X"2C",X"20",X"01",
		X"90",X"4C",X"10",X"01",X"20",X"1C",X"60",X"3C",X"20",X"01",X"20",X"2C",X"40",X"2C",X"2C",X"20",
		X"01",X"20",X"3C",X"20",X"4C",X"30",X"01",X"10",X"5C",X"20",X"3C",X"30",X"01",X"10",X"3C",X"10",
		X"24",X"4C",X"30",X"01",X"10",X"3C",X"54",X"24",X"30",X"01",X"40",X"64",X"40",X"01",X"60",X"2C",
		X"00",X"70",X"01",X"70",X"01",X"70",X"01",X"20",X"37",X"20",X"01",X"10",X"57",X"10",X"01",X"77",
		X"01",X"27",X"4C",X"17",X"01",X"37",X"2C",X"27",X"01",X"10",X"57",X"10",X"00",X"01",X"01",X"01",
		X"01",X"E0",X"01",X"E0",X"01",X"E0",X"01",X"E0",X"01",X"30",X"2E",X"30",X"2E",X"40",X"01",X"40",
		X"4E",X"60",X"01",X"20",X"8E",X"40",X"01",X"10",X"4E",X"4C",X"2E",X"30",X"01",X"10",X"3E",X"2C",
		X"24",X"2C",X"1E",X"30",X"01",X"10",X"5E",X"2C",X"3E",X"30",X"01",X"60",X"2C",X"00",X"01",X"01",
		X"01",X"70",X"01",X"70",X"01",X"70",X"01",X"20",X"3E",X"20",X"01",X"10",X"5E",X"10",X"01",X"3E",
		X"2C",X"2E",X"01",X"10",X"5E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"38",X"D8",X"7E",X"39",X"DA",X"7E",X"3C",X"B2",X"7E",X"3C",X"AC",X"7E",X"3C",X"58",X"7E",
		X"3C",X"7D",X"7E",X"3C",X"8E",X"7E",X"3C",X"8C",X"7E",X"3C",X"96",X"7E",X"3C",X"A4",X"7E",X"3C",
		X"A2",X"7E",X"3C",X"EB",X"7E",X"3E",X"CE",X"7E",X"3E",X"C8",X"7E",X"3E",X"C2",X"7E",X"3F",X"49",
		X"7E",X"3F",X"5E",X"7E",X"40",X"86",X"7E",X"42",X"16",X"7E",X"3B",X"5D",X"7E",X"39",X"92",X"7E",
		X"3A",X"08",X"7E",X"39",X"9F",X"7E",X"39",X"5D",X"7E",X"39",X"C5",X"7E",X"38",X"6B",X"7D",X"BF",
		X"35",X"27",X"3E",X"86",X"04",X"BD",X"5D",X"9F",X"BD",X"37",X"BC",X"8E",X"26",X"20",X"86",X"58",
		X"C6",X"11",X"BD",X"46",X"23",X"8E",X"14",X"CA",X"86",X"5A",X"C6",X"99",X"BD",X"46",X"2C",X"BE",
		X"5D",X"A5",X"BD",X"5D",X"90",X"6F",X"C8",X"32",X"86",X"1E",X"BD",X"5D",X"9F",X"7F",X"98",X"68",
		X"6A",X"C8",X"32",X"27",X"0F",X"AE",X"C4",X"A6",X"05",X"81",X"41",X"27",X"EB",X"81",X"42",X"27",
		X"E7",X"7E",X"5D",X"93",X"86",X"42",X"BD",X"5D",X"A2",X"86",X"03",X"BD",X"5D",X"9F",X"20",X"F1",
		X"34",X"02",X"A6",X"80",X"1E",X"12",X"BD",X"3C",X"96",X"1E",X"12",X"5A",X"26",X"F4",X"35",X"82",
		X"8E",X"CC",X"00",X"6F",X"80",X"8C",X"D0",X"00",X"26",X"F9",X"39",X"34",X"36",X"8E",X"38",X"92",
		X"10",X"8E",X"CC",X"00",X"C6",X"12",X"8D",X"D8",X"35",X"B6",X"34",X"36",X"8E",X"38",X"A4",X"10",
		X"8E",X"CC",X"24",X"C6",X"34",X"8D",X"C9",X"BD",X"39",X"76",X"8E",X"CC",X"8E",X"BD",X"3C",X"96",
		X"35",X"B6",X"30",X"03",X"25",X"03",X"01",X"04",X"01",X"01",X"00",X"00",X"05",X"03",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"1A",X"1C",X"0F",X"1D",X"0F",
		X"18",X"1E",X"0F",X"0E",X"0A",X"0C",X"23",X"2C",X"0A",X"0A",X"0A",X"0A",X"0A",X"21",X"13",X"16",
		X"16",X"13",X"0B",X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",
		X"1D",X"0A",X"13",X"18",X"0D",X"2D",X"25",X"29",X"BD",X"39",X"5D",X"BD",X"3C",X"58",X"B6",X"C8",
		X"0C",X"85",X"02",X"26",X"F9",X"B6",X"CC",X"1B",X"84",X"0F",X"27",X"11",X"7F",X"CC",X"1B",X"BD",
		X"39",X"5D",X"BD",X"3C",X"58",X"BD",X"39",X"B5",X"86",X"40",X"BD",X"F0",X"09",X"B6",X"CC",X"1D",
		X"84",X"0F",X"27",X"0D",X"7F",X"CC",X"1D",X"8D",X"54",X"BD",X"3A",X"28",X"86",X"40",X"BD",X"F0",
		X"09",X"B6",X"CC",X"21",X"84",X"0F",X"27",X"1E",X"7F",X"CC",X"21",X"8D",X"40",X"BD",X"3C",X"58",
		X"86",X"0A",X"BD",X"46",X"32",X"BD",X"41",X"10",X"96",X"20",X"BD",X"F0",X"09",X"BD",X"39",X"76",
		X"8E",X"CC",X"8E",X"BD",X"3C",X"96",X"B6",X"CC",X"1F",X"84",X"0F",X"27",X"0A",X"7F",X"CC",X"1F",
		X"8D",X"1B",X"8D",X"08",X"7E",X"F0",X"06",X"8D",X"03",X"7E",X"F0",X"0F",X"B6",X"CC",X"19",X"84",
		X"0F",X"27",X"09",X"7C",X"CC",X"8C",X"7C",X"CC",X"8C",X"7F",X"CC",X"19",X"39",X"34",X"12",X"8D",
		X"08",X"8E",X"CC",X"8C",X"BD",X"3C",X"96",X"35",X"92",X"34",X"34",X"8E",X"CC",X"00",X"10",X"8E",
		X"CC",X"24",X"8D",X"09",X"35",X"B4",X"8E",X"CC",X"24",X"10",X"8E",X"CC",X"8C",X"10",X"BF",X"BF",
		X"15",X"4F",X"E6",X"80",X"C4",X"0F",X"34",X"04",X"AB",X"E0",X"BC",X"BF",X"15",X"26",X"F3",X"8B",
		X"37",X"39",X"8D",X"D5",X"34",X"02",X"8E",X"CC",X"8C",X"BD",X"3C",X"7D",X"A1",X"E0",X"39",X"8E",
		X"CD",X"02",X"C6",X"04",X"A6",X"80",X"84",X"0F",X"81",X"09",X"23",X"03",X"5A",X"27",X"06",X"8C",
		X"CD",X"3E",X"26",X"F0",X"39",X"86",X"0D",X"BD",X"46",X"32",X"8E",X"CD",X"02",X"6F",X"80",X"8C",
		X"CD",X"3E",X"26",X"F9",X"39",X"8D",X"05",X"27",X"FB",X"7E",X"38",X"7A",X"BD",X"39",X"76",X"34",
		X"02",X"8E",X"CC",X"8E",X"BD",X"3C",X"7D",X"A1",X"E0",X"39",X"86",X"18",X"B7",X"BF",X"22",X"86",
		X"3F",X"B7",X"C8",X"0E",X"86",X"08",X"BD",X"F0",X"09",X"B6",X"C8",X"0C",X"85",X"08",X"27",X"17",
		X"7A",X"BF",X"22",X"26",X"EF",X"10",X"8E",X"CD",X"3E",X"8E",X"3A",X"82",X"C6",X"17",X"BD",X"38",
		X"50",X"BD",X"3B",X"24",X"7F",X"C8",X"0E",X"39",X"10",X"8E",X"CD",X"74",X"C6",X"08",X"BD",X"3B",
		X"4B",X"A8",X"26",X"84",X"0F",X"27",X"03",X"5A",X"27",X"0E",X"86",X"39",X"B7",X"CB",X"FF",X"31",
		X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"E7",X"39",X"86",X"39",X"B7",X"CB",X"FF",X"10",X"8E",X"3A",
		X"82",X"8E",X"CD",X"3E",X"C6",X"14",X"A6",X"A0",X"BD",X"3C",X"96",X"5A",X"26",X"F8",X"C6",X"29",
		X"8D",X"1C",X"BD",X"3B",X"24",X"10",X"8E",X"CD",X"74",X"BD",X"3B",X"43",X"86",X"39",X"B7",X"CB",
		X"FF",X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"F0",X"86",X"0E",X"7E",X"46",X"32",X"E7",X"E2",
		X"A6",X"A0",X"BD",X"3C",X"96",X"A6",X"A0",X"BD",X"3C",X"96",X"A6",X"A0",X"BD",X"3C",X"96",X"4F",
		X"5F",X"ED",X"84",X"ED",X"04",X"ED",X"06",X"5C",X"ED",X"02",X"30",X"08",X"6A",X"E4",X"26",X"E0",
		X"35",X"84",X"1D",X"1A",X"16",X"0B",X"1E",X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",
		X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"21",X"13",X"16",X"17",X"1C",X"1D",X"14",X"1C",X"18",X"12",
		X"0F",X"0D",X"17",X"0C",X"1D",X"1A",X"10",X"24",X"14",X"13",X"16",X"0D",X"21",X"15",X"1C",X"1D",
		X"17",X"0F",X"0A",X"24",X"15",X"0F",X"18",X"20",X"1D",X"17",X"0D",X"1C",X"0C",X"1A",X"20",X"0B",
		X"11",X"21",X"21",X"1C",X"19",X"18",X"14",X"19",X"0F",X"1E",X"13",X"17",X"1C",X"1D",X"17",X"14",
		X"13",X"17",X"20",X"13",X"0D",X"16",X"0F",X"19",X"0C",X"1F",X"24",X"14",X"14",X"15",X"1C",X"0F",
		X"18",X"18",X"0A",X"10",X"14",X"1C",X"18",X"12",X"0F",X"0D",X"17",X"0C",X"1D",X"1A",X"10",X"24",
		X"14",X"13",X"16",X"1C",X"20",X"1E",X"15",X"0B",X"23",X"14",X"11",X"16",X"1C",X"0B",X"17",X"12",
		X"0F",X"0D",X"15",X"20",X"0E",X"0F",X"14",X"1D",X"20",X"0B",X"22",X"0E",X"1C",X"14",X"14",X"0B",
		X"23",X"12",X"17",X"0C",X"00",X"00",X"40",X"00",X"34",X"34",X"8E",X"3B",X"11",X"C6",X"07",X"BD",
		X"38",X"50",X"35",X"B4",X"34",X"02",X"8D",X"05",X"B7",X"CD",X"6C",X"35",X"82",X"34",X"10",X"8E",
		X"CD",X"3E",X"4F",X"AB",X"84",X"30",X"01",X"8C",X"CD",X"6C",X"27",X"F9",X"8C",X"CD",X"74",X"26",
		X"F2",X"35",X"90",X"34",X"02",X"8D",X"04",X"A7",X"26",X"35",X"82",X"34",X"24",X"C6",X"0E",X"4F",
		X"C1",X"08",X"27",X"02",X"AB",X"A4",X"31",X"21",X"5A",X"26",X"F5",X"35",X"A4",X"86",X"32",X"34",
		X"02",X"10",X"8E",X"CD",X"74",X"8D",X"E4",X"A8",X"26",X"84",X"0F",X"27",X"0F",X"BD",X"3C",X"2D",
		X"7F",X"CD",X"00",X"7F",X"CD",X"01",X"6A",X"E4",X"27",X"12",X"20",X"E9",X"86",X"03",X"C6",X"04",
		X"8D",X"65",X"25",X"E9",X"31",X"2E",X"10",X"8C",X"CF",X"A4",X"25",X"D9",X"35",X"02",X"10",X"8E",
		X"3A",X"9C",X"8E",X"CF",X"A4",X"C6",X"06",X"BD",X"3A",X"5E",X"8D",X"91",X"B8",X"CD",X"6C",X"84",
		X"0F",X"27",X"02",X"8D",X"0F",X"10",X"8E",X"CD",X"3E",X"86",X"17",X"C6",X"04",X"8D",X"38",X"24",
		X"02",X"8D",X"01",X"39",X"8E",X"CD",X"3E",X"86",X"0A",X"BD",X"3C",X"96",X"8C",X"CD",X"66",X"25",
		X"F8",X"8E",X"CD",X"74",X"10",X"8E",X"CD",X"3E",X"86",X"06",X"BD",X"3C",X"4D",X"10",X"8E",X"CD",
		X"66",X"8D",X"7A",X"8E",X"CD",X"7A",X"10",X"8E",X"CD",X"6C",X"86",X"08",X"8D",X"6F",X"BD",X"3B",
		X"24",X"10",X"8E",X"CD",X"74",X"20",X"46",X"34",X"16",X"C6",X"39",X"F7",X"CB",X"FF",X"1F",X"21",
		X"BD",X"3C",X"8E",X"C1",X"0A",X"25",X"32",X"C1",X"24",X"22",X"2E",X"4A",X"26",X"F2",X"A6",X"61",
		X"BD",X"3C",X"8E",X"C4",X"0F",X"C1",X"09",X"22",X"20",X"4A",X"BD",X"3C",X"8E",X"34",X"04",X"C4",
		X"0F",X"C1",X"09",X"35",X"04",X"22",X"12",X"C4",X"F0",X"C1",X"99",X"22",X"0C",X"4A",X"26",X"EA",
		X"1C",X"FE",X"86",X"39",X"B7",X"CB",X"FF",X"35",X"96",X"1A",X"01",X"20",X"F5",X"34",X"36",X"30",
		X"2E",X"8C",X"CF",X"A4",X"24",X"0F",X"86",X"0E",X"8D",X"13",X"31",X"2E",X"30",X"0E",X"86",X"39",
		X"B7",X"CB",X"FF",X"20",X"EC",X"BD",X"3B",X"18",X"BD",X"3B",X"43",X"35",X"B6",X"34",X"36",X"E6",
		X"80",X"E7",X"A0",X"4A",X"26",X"F9",X"35",X"B6",X"34",X"76",X"CC",X"00",X"00",X"1F",X"01",X"1F",
		X"02",X"CE",X"98",X"00",X"86",X"39",X"36",X"34",X"36",X"34",X"36",X"34",X"36",X"34",X"36",X"34",
		X"36",X"34",X"B7",X"CB",X"FF",X"11",X"83",X"98",X"00",X"25",X"EB",X"35",X"F6",X"A6",X"01",X"84",
		X"0F",X"34",X"02",X"A6",X"81",X"48",X"48",X"48",X"48",X"AB",X"E0",X"39",X"8D",X"EF",X"34",X"02",
		X"8D",X"EB",X"1F",X"89",X"35",X"82",X"34",X"02",X"A7",X"01",X"44",X"44",X"44",X"44",X"A7",X"81",
		X"35",X"82",X"8D",X"F2",X"34",X"02",X"1F",X"98",X"8D",X"EC",X"35",X"82",X"34",X"16",X"86",X"01",
		X"20",X"02",X"34",X"16",X"C4",X"0F",X"58",X"34",X"04",X"58",X"EB",X"E0",X"8E",X"CC",X"FC",X"3A",
		X"8D",X"CC",X"34",X"04",X"8D",X"C8",X"34",X"04",X"8D",X"C4",X"34",X"04",X"AB",X"E4",X"19",X"A7",
		X"E4",X"A6",X"61",X"89",X"00",X"19",X"A7",X"61",X"A6",X"62",X"89",X"00",X"19",X"30",X"1A",X"8D",
		X"B5",X"35",X"04",X"35",X"02",X"8D",X"BB",X"35",X"02",X"35",X"96",X"86",X"0F",X"BD",X"46",X"32",
		X"7F",X"BF",X"15",X"8E",X"11",X"70",X"CC",X"F1",X"22",X"10",X"8E",X"CD",X"3E",X"10",X"BC",X"BF",
		X"2A",X"26",X"04",X"C6",X"44",X"20",X"08",X"10",X"BC",X"BF",X"2E",X"26",X"02",X"C6",X"55",X"BD",
		X"46",X"26",X"86",X"2A",X"BD",X"46",X"20",X"30",X"89",X"03",X"00",X"86",X"15",X"B7",X"BF",X"1C",
		X"7A",X"BF",X"1C",X"27",X"1E",X"1E",X"12",X"BD",X"37",X"BF",X"81",X"0A",X"2E",X"0B",X"7D",X"BF",
		X"15",X"26",X"09",X"10",X"BF",X"BF",X"15",X"20",X"03",X"7F",X"BF",X"15",X"1E",X"12",X"BD",X"46",
		X"20",X"20",X"DD",X"7D",X"BF",X"15",X"27",X"03",X"BE",X"BF",X"15",X"86",X"04",X"B7",X"BF",X"1C",
		X"10",X"8E",X"CD",X"6C",X"1E",X"12",X"BD",X"37",X"BF",X"1E",X"12",X"8A",X"F0",X"85",X"0F",X"26",
		X"02",X"8A",X"0F",X"BD",X"46",X"26",X"7A",X"BF",X"1C",X"1E",X"12",X"BD",X"37",X"BF",X"1E",X"12",
		X"BD",X"46",X"26",X"7A",X"BF",X"1C",X"26",X"F1",X"8E",X"13",X"80",X"C6",X"33",X"CE",X"46",X"2F",
		X"FF",X"BF",X"1F",X"CE",X"46",X"29",X"86",X"0D",X"B7",X"BF",X"1C",X"86",X"02",X"B7",X"BF",X"22",
		X"86",X"07",X"B7",X"BF",X"21",X"86",X"0F",X"B7",X"BF",X"27",X"8D",X"53",X"8E",X"3D",X"80",X"86",
		X"0D",X"B7",X"BF",X"1C",X"86",X"15",X"B7",X"BF",X"22",X"8D",X"44",X"8E",X"67",X"80",X"86",X"0D",
		X"B7",X"BF",X"1C",X"86",X"28",X"B7",X"BF",X"22",X"8D",X"35",X"8E",X"13",X"36",X"10",X"8E",X"CF",
		X"A4",X"C6",X"11",X"CE",X"46",X"26",X"FF",X"BF",X"1F",X"CE",X"46",X"20",X"86",X"03",X"B7",X"BF",
		X"1C",X"86",X"01",X"B7",X"BF",X"22",X"86",X"0A",X"B7",X"BF",X"21",X"86",X"15",X"B7",X"BF",X"27",
		X"8D",X"0D",X"8E",X"53",X"36",X"86",X"03",X"B7",X"BF",X"1C",X"86",X"04",X"B7",X"BF",X"22",X"BF",
		X"BF",X"19",X"34",X"04",X"C6",X"03",X"F7",X"BF",X"29",X"5C",X"F7",X"BF",X"26",X"E6",X"E4",X"10",
		X"BC",X"BF",X"2A",X"27",X"06",X"10",X"BC",X"BF",X"2C",X"26",X"02",X"C6",X"44",X"10",X"BC",X"BF",
		X"2E",X"27",X"06",X"10",X"BC",X"BF",X"30",X"26",X"02",X"C6",X"55",X"B6",X"BF",X"22",X"85",X"F0",
		X"26",X"02",X"8A",X"F0",X"AD",X"9F",X"BF",X"1F",X"86",X"2A",X"AD",X"C4",X"86",X"0A",X"AD",X"C4",
		X"1E",X"12",X"BD",X"37",X"BF",X"1E",X"12",X"AD",X"C4",X"7A",X"BF",X"29",X"26",X"F2",X"BF",X"BF",
		X"15",X"BE",X"BF",X"19",X"1E",X"01",X"F6",X"BF",X"16",X"BB",X"BF",X"27",X"1E",X"01",X"7F",X"BF",
		X"1D",X"1E",X"12",X"BD",X"37",X"BF",X"1E",X"12",X"7D",X"BF",X"1D",X"26",X"1B",X"34",X"02",X"86",
		X"04",X"B1",X"BF",X"26",X"26",X"04",X"35",X"02",X"20",X"06",X"35",X"02",X"85",X"F0",X"26",X"08",
		X"8A",X"F0",X"85",X"0F",X"26",X"02",X"8A",X"0F",X"B7",X"BF",X"1D",X"73",X"BF",X"1D",X"AD",X"9F",
		X"BF",X"1F",X"7A",X"BF",X"26",X"26",X"CA",X"BF",X"BF",X"15",X"BE",X"BF",X"19",X"1E",X"01",X"F6",
		X"BF",X"16",X"FB",X"BF",X"21",X"1E",X"01",X"B6",X"BF",X"22",X"8B",X"01",X"19",X"B7",X"BF",X"22",
		X"7A",X"BF",X"1C",X"35",X"04",X"10",X"26",X"FF",X"49",X"39",X"34",X"12",X"BB",X"BF",X"32",X"19",
		X"24",X"02",X"86",X"99",X"B7",X"BF",X"32",X"8E",X"CD",X"00",X"BD",X"3C",X"96",X"35",X"12",X"7E",
		X"5D",X"96",X"34",X"16",X"C6",X"03",X"20",X"0A",X"34",X"16",X"C6",X"02",X"20",X"04",X"34",X"16",
		X"C6",X"01",X"BD",X"3C",X"AC",X"58",X"8E",X"CC",X"06",X"3A",X"BD",X"3C",X"8E",X"8D",X"6A",X"B6",
		X"BF",X"34",X"34",X"04",X"AB",X"E4",X"B7",X"BF",X"34",X"B6",X"BF",X"33",X"AB",X"E0",X"B7",X"BF",
		X"33",X"8E",X"CC",X"12",X"BD",X"3C",X"8E",X"8D",X"50",X"34",X"04",X"A1",X"E0",X"24",X"02",X"35",
		X"96",X"8E",X"CC",X"0E",X"BD",X"3C",X"8E",X"8D",X"40",X"8D",X"28",X"34",X"02",X"F7",X"BF",X"33",
		X"8E",X"CC",X"10",X"BD",X"3C",X"8E",X"B6",X"BF",X"34",X"8D",X"2E",X"8D",X"16",X"4D",X"27",X"06",
		X"7F",X"BF",X"33",X"7F",X"BF",X"34",X"AB",X"E0",X"19",X"C6",X"04",X"BD",X"3C",X"B2",X"BD",X"3E",
		X"AA",X"35",X"96",X"34",X"04",X"5D",X"26",X"03",X"4F",X"35",X"84",X"1E",X"89",X"86",X"99",X"8B",
		X"01",X"19",X"E0",X"E4",X"24",X"F9",X"EB",X"E0",X"39",X"34",X"02",X"4F",X"C1",X"10",X"25",X"06",
		X"8B",X"0A",X"C0",X"10",X"20",X"F6",X"34",X"04",X"AB",X"E0",X"1F",X"89",X"35",X"82",X"34",X"04",
		X"1F",X"89",X"4F",X"C1",X"0A",X"25",X"07",X"8B",X"10",X"19",X"C0",X"0A",X"20",X"F5",X"34",X"04",
		X"AB",X"E0",X"19",X"35",X"84",X"4F",X"E6",X"21",X"27",X"11",X"34",X"04",X"CB",X"0E",X"E6",X"A5",
		X"58",X"BE",X"46",X"38",X"AB",X"95",X"35",X"04",X"5A",X"26",X"EF",X"AE",X"28",X"30",X"8B",X"AF",
		X"2A",X"C6",X"0F",X"EB",X"21",X"A6",X"A5",X"BD",X"40",X"35",X"E6",X"24",X"F7",X"C8",X"07",X"F6",
		X"C8",X"04",X"C4",X"43",X"26",X"08",X"E6",X"2E",X"27",X"70",X"6A",X"2E",X"20",X"6C",X"8E",X"3F",
		X"B6",X"AF",X"26",X"1C",X"FE",X"39",X"34",X"04",X"E6",X"24",X"F7",X"C8",X"07",X"F6",X"C8",X"04",
		X"C4",X"43",X"E1",X"E4",X"35",X"04",X"26",X"52",X"C5",X"FD",X"26",X"0D",X"8D",X"5F",X"A1",X"22",
		X"26",X"04",X"A6",X"23",X"20",X"12",X"4A",X"20",X"0F",X"C5",X"40",X"26",X"13",X"8D",X"4E",X"A1",
		X"23",X"26",X"04",X"A6",X"22",X"20",X"01",X"4C",X"E6",X"2E",X"27",X"2E",X"6A",X"2E",X"20",X"2A",
		X"E6",X"2E",X"26",X"F8",X"C6",X"02",X"E7",X"2E",X"81",X"25",X"26",X"0E",X"6D",X"21",X"27",X"1A",
		X"8D",X"2B",X"8D",X"2C",X"6C",X"A4",X"6A",X"21",X"20",X"12",X"8D",X"24",X"6C",X"21",X"6A",X"A4",
		X"26",X"08",X"1A",X"01",X"8E",X"3F",X"75",X"AF",X"26",X"39",X"8D",X"04",X"1C",X"FE",X"20",X"F4",
		X"C6",X"0F",X"EB",X"21",X"A7",X"A5",X"E6",X"25",X"AE",X"2A",X"7E",X"46",X"20",X"5F",X"20",X"F8",
		X"34",X"27",X"5F",X"20",X"04",X"34",X"27",X"E6",X"25",X"1A",X"F0",X"F7",X"CA",X"01",X"CC",X"40",
		X"75",X"FD",X"CA",X"02",X"AE",X"2A",X"30",X"08",X"CC",X"04",X"02",X"8D",X"19",X"CC",X"40",X"76",
		X"FD",X"CA",X"02",X"E6",X"A4",X"5A",X"2F",X"0C",X"4F",X"1F",X"02",X"CC",X"03",X"01",X"8D",X"06",
		X"31",X"3F",X"26",X"F7",X"35",X"A7",X"FD",X"CA",X"06",X"BF",X"CA",X"04",X"C6",X"1A",X"F7",X"CA",
		X"00",X"5F",X"30",X"8B",X"39",X"11",X"11",X"11",X"10",X"11",X"11",X"11",X"10",X"34",X"06",X"86",
		X"04",X"BD",X"F0",X"09",X"35",X"86",X"C6",X"66",X"F7",X"BF",X"29",X"C6",X"88",X"8D",X"04",X"C6",
		X"9A",X"20",X"21",X"34",X"36",X"8E",X"CC",X"88",X"BD",X"37",X"BF",X"1F",X"02",X"8E",X"CC",X"24",
		X"F6",X"BF",X"29",X"BD",X"37",X"BF",X"1E",X"12",X"BD",X"46",X"20",X"1E",X"12",X"8C",X"CC",X"56",
		X"26",X"F1",X"35",X"B6",X"34",X"36",X"8E",X"CC",X"8A",X"BD",X"37",X"BF",X"1F",X"02",X"8E",X"CC",
		X"56",X"F6",X"BF",X"29",X"BD",X"37",X"BF",X"1E",X"12",X"BD",X"46",X"20",X"1E",X"12",X"8C",X"CC",
		X"88",X"26",X"F1",X"35",X"B6",X"10",X"8E",X"B0",X"00",X"AF",X"28",X"CC",X"3F",X"75",X"ED",X"26",
		X"C6",X"02",X"E7",X"2E",X"C6",X"19",X"E7",X"A4",X"C6",X"14",X"86",X"0A",X"30",X"2F",X"A7",X"80",
		X"5A",X"26",X"FB",X"E7",X"21",X"E7",X"22",X"6F",X"2F",X"86",X"31",X"A7",X"23",X"86",X"3C",X"A7",
		X"24",X"86",X"77",X"A7",X"25",X"AD",X"B8",X"06",X"25",X"05",X"BD",X"40",X"7D",X"20",X"F6",X"39",
		X"8E",X"25",X"60",X"8D",X"C0",X"C6",X"19",X"8E",X"CC",X"24",X"31",X"2F",X"A6",X"A0",X"BD",X"3C",
		X"96",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",X"88",X"BD",X"3C",X"96",X"C6",X"88",X"8D",X"34",
		X"86",X"31",X"C6",X"22",X"8E",X"48",X"6A",X"BD",X"46",X"20",X"CE",X"41",X"74",X"8E",X"CC",X"88",
		X"BD",X"3C",X"8E",X"BD",X"41",X"D5",X"F7",X"BF",X"37",X"7F",X"BF",X"29",X"C6",X"60",X"BD",X"40",
		X"93",X"B6",X"BF",X"37",X"8E",X"CC",X"88",X"BD",X"3C",X"96",X"86",X"22",X"B7",X"BF",X"29",X"BD",
		X"40",X"93",X"20",X"D9",X"86",X"51",X"8E",X"25",X"90",X"BD",X"46",X"23",X"86",X"52",X"8E",X"25",
		X"A0",X"7E",X"46",X"23",X"86",X"31",X"C6",X"00",X"8E",X"48",X"6A",X"BD",X"46",X"20",X"8D",X"E4",
		X"8E",X"25",X"70",X"BD",X"40",X"D5",X"C6",X"19",X"8E",X"CC",X"56",X"31",X"2F",X"A6",X"A0",X"BD",
		X"3C",X"96",X"5A",X"26",X"F8",X"86",X"25",X"8E",X"CC",X"8A",X"BD",X"3C",X"96",X"C6",X"88",X"8D",
		X"C3",X"86",X"31",X"C6",X"22",X"8E",X"48",X"7A",X"BD",X"46",X"20",X"CE",X"41",X"D4",X"8E",X"CC",
		X"8A",X"BD",X"3C",X"8E",X"8D",X"1F",X"F7",X"BF",X"37",X"7F",X"BF",X"29",X"C6",X"70",X"BD",X"40",
		X"B4",X"B6",X"BF",X"37",X"8E",X"CC",X"8A",X"BD",X"3C",X"96",X"86",X"22",X"B7",X"BF",X"29",X"BD",
		X"40",X"B4",X"20",X"DA",X"39",X"B6",X"C8",X"0C",X"85",X"02",X"27",X"04",X"32",X"62",X"6E",X"C4",
		X"B6",X"C8",X"04",X"84",X"03",X"BD",X"40",X"7D",X"34",X"02",X"B6",X"C8",X"04",X"84",X"03",X"A1",
		X"E4",X"35",X"02",X"26",X"E0",X"4D",X"27",X"DD",X"85",X"FE",X"26",X"06",X"C1",X"18",X"27",X"D5",
		X"5A",X"39",X"C1",X"40",X"27",X"CF",X"5C",X"39",X"A6",X"84",X"84",X"F0",X"27",X"07",X"CC",X"99",
		X"99",X"ED",X"81",X"ED",X"81",X"39",X"7F",X"BF",X"35",X"B6",X"CC",X"23",X"44",X"25",X"03",X"7E",
		X"5D",X"93",X"8E",X"99",X"0C",X"8D",X"E1",X"8E",X"99",X"15",X"8D",X"DC",X"7D",X"98",X"23",X"27",
		X"5C",X"8E",X"99",X"0C",X"10",X"8E",X"99",X"15",X"BD",X"45",X"73",X"25",X"50",X"1E",X"21",X"BD",
		X"45",X"37",X"24",X"24",X"7C",X"BF",X"35",X"8E",X"44",X"C1",X"86",X"42",X"BD",X"5D",X"99",X"1F",
		X"12",X"86",X"10",X"A7",X"24",X"86",X"01",X"A7",X"A8",X"31",X"8E",X"99",X"15",X"AF",X"A8",X"2D",
		X"8E",X"70",X"A0",X"AF",X"A8",X"2F",X"20",X"12",X"8E",X"99",X"15",X"AF",X"C8",X"2D",X"8E",X"70",
		X"A0",X"AF",X"C8",X"2F",X"86",X"01",X"C6",X"42",X"8D",X"69",X"8E",X"99",X"0C",X"AF",X"C8",X"2D",
		X"8E",X"20",X"A0",X"AF",X"C8",X"2F",X"4F",X"C6",X"41",X"8D",X"58",X"20",X"53",X"8E",X"99",X"0C",
		X"BD",X"45",X"37",X"24",X"23",X"7C",X"BF",X"35",X"8E",X"44",X"C1",X"86",X"42",X"BD",X"5D",X"99",
		X"1F",X"12",X"86",X"10",X"A7",X"24",X"4F",X"A7",X"A8",X"31",X"8E",X"99",X"0C",X"AF",X"A8",X"2D",
		X"8E",X"20",X"A0",X"AF",X"A8",X"2F",X"20",X"11",X"8E",X"99",X"0C",X"AF",X"C8",X"2D",X"8E",X"20",
		X"A0",X"AF",X"C8",X"2F",X"4F",X"C6",X"42",X"8D",X"1A",X"7D",X"98",X"23",X"27",X"12",X"8E",X"99",
		X"15",X"AF",X"C8",X"2D",X"8E",X"70",X"A0",X"AF",X"C8",X"2F",X"86",X"01",X"C6",X"41",X"8D",X"03",
		X"7E",X"37",X"FE",X"BD",X"45",X"3D",X"24",X"26",X"7C",X"BF",X"35",X"34",X"02",X"8E",X"43",X"39",
		X"1F",X"98",X"5F",X"BD",X"5D",X"99",X"1F",X"12",X"86",X"10",X"A7",X"24",X"35",X"02",X"A7",X"A8",
		X"31",X"AE",X"C8",X"2D",X"AF",X"A8",X"2D",X"AE",X"C8",X"2F",X"AF",X"A8",X"2F",X"39",X"BD",X"45",
		X"5A",X"24",X"25",X"7C",X"BF",X"35",X"34",X"02",X"8E",X"43",X"39",X"1F",X"98",X"5F",X"BD",X"5D",
		X"99",X"1F",X"12",X"86",X"08",X"A7",X"24",X"35",X"02",X"A7",X"A8",X"31",X"AE",X"C8",X"2D",X"AF",
		X"A8",X"2D",X"AE",X"C8",X"2F",X"AF",X"A8",X"2F",X"39",X"6F",X"C8",X"2C",X"E6",X"C8",X"31",X"26",
		X"0B",X"8E",X"0A",X"B0",X"C6",X"3C",X"34",X"04",X"C6",X"44",X"20",X"09",X"8E",X"58",X"B0",X"C6",
		X"34",X"34",X"04",X"C6",X"55",X"86",X"57",X"BD",X"46",X"23",X"1F",X"98",X"31",X"47",X"35",X"04",
		X"E7",X"24",X"8E",X"43",X"6D",X"AF",X"2C",X"AE",X"C8",X"2F",X"7E",X"45",X"AC",X"A6",X"45",X"81",
		X"42",X"27",X"21",X"ED",X"C8",X"32",X"AF",X"C8",X"34",X"10",X"AF",X"C8",X"36",X"86",X"01",X"BD",
		X"5D",X"9F",X"AE",X"C4",X"A6",X"05",X"81",X"42",X"27",X"F3",X"EC",X"C8",X"32",X"AE",X"C8",X"34",
		X"10",X"AE",X"C8",X"36",X"BD",X"45",X"3D",X"24",X"15",X"6D",X"C8",X"31",X"26",X"06",X"10",X"BF",
		X"BF",X"2C",X"20",X"04",X"10",X"BF",X"BF",X"30",X"8E",X"CF",X"EA",X"BD",X"44",X"90",X"BD",X"45",
		X"5A",X"24",X"19",X"6D",X"C8",X"2C",X"27",X"1D",X"30",X"47",X"30",X"0F",X"10",X"8E",X"CD",X"66",
		X"C6",X"03",X"BD",X"38",X"50",X"BD",X"3B",X"24",X"86",X"05",X"8D",X"79",X"24",X"74",X"1F",X"12",
		X"BD",X"3C",X"2D",X"20",X"55",X"30",X"A9",X"32",X"9A",X"26",X"2E",X"8E",X"CF",X"96",X"BD",X"44",
		X"AB",X"31",X"26",X"AE",X"C8",X"2D",X"C6",X"04",X"BD",X"38",X"50",X"10",X"8E",X"CD",X"3E",X"6D",
		X"C8",X"31",X"26",X"06",X"10",X"BF",X"BF",X"2A",X"20",X"04",X"10",X"BF",X"BF",X"2E",X"30",X"47",
		X"30",X"0F",X"C6",X"14",X"BD",X"38",X"50",X"20",X"AF",X"BD",X"44",X"49",X"34",X"01",X"34",X"10",
		X"10",X"AC",X"E1",X"22",X"11",X"8D",X"79",X"6D",X"C8",X"31",X"26",X"06",X"10",X"BF",X"BF",X"2A",
		X"20",X"04",X"10",X"BF",X"BF",X"2E",X"35",X"01",X"24",X"18",X"8E",X"BF",X"2A",X"31",X"47",X"AE",
		X"C8",X"2F",X"30",X"89",X"EA",X"F6",X"86",X"59",X"E6",X"25",X"BD",X"46",X"23",X"86",X"60",X"BD",
		X"5D",X"9F",X"7E",X"5D",X"9C",X"34",X"26",X"20",X"0C",X"34",X"26",X"8E",X"CD",X"66",X"8D",X"26",
		X"86",X"04",X"25",X"01",X"4C",X"B7",X"BF",X"15",X"8E",X"CD",X"74",X"8D",X"19",X"24",X"05",X"7A",
		X"BF",X"15",X"27",X"0E",X"30",X"0E",X"8C",X"CF",X"A4",X"25",X"F0",X"8E",X"CF",X"96",X"1C",X"FE",
		X"35",X"A6",X"1A",X"01",X"35",X"A6",X"34",X"10",X"31",X"47",X"31",X"2F",X"C6",X"03",X"BD",X"3C",
		X"7D",X"A1",X"A0",X"26",X"07",X"5A",X"26",X"F6",X"1A",X"01",X"35",X"90",X"1C",X"FE",X"35",X"90",
		X"34",X"20",X"BD",X"44",X"AB",X"30",X"47",X"30",X"0F",X"C6",X"03",X"BD",X"38",X"50",X"AE",X"C8",
		X"2D",X"C6",X"04",X"BD",X"38",X"50",X"35",X"20",X"7E",X"3B",X"43",X"34",X"30",X"1F",X"12",X"10",
		X"AC",X"62",X"27",X"0B",X"30",X"32",X"86",X"0E",X"BD",X"3C",X"4D",X"31",X"32",X"20",X"F0",X"35",
		X"B0",X"6C",X"C8",X"2C",X"31",X"47",X"A6",X"C8",X"31",X"26",X"08",X"86",X"3C",X"A7",X"24",X"86",
		X"44",X"20",X"06",X"86",X"34",X"A7",X"24",X"86",X"55",X"1F",X"89",X"86",X"56",X"8E",X"1E",X"5B",
		X"BD",X"46",X"23",X"1F",X"98",X"8E",X"44",X"ED",X"AF",X"2C",X"7E",X"45",X"9E",X"30",X"2F",X"10",
		X"8E",X"CD",X"3E",X"C6",X"14",X"BD",X"38",X"50",X"10",X"8E",X"CD",X"66",X"8E",X"CF",X"96",X"BD",
		X"44",X"AB",X"10",X"8E",X"CD",X"74",X"BD",X"3B",X"43",X"AE",X"C8",X"2D",X"10",X"8E",X"CD",X"6C",
		X"C6",X"04",X"BD",X"38",X"50",X"8E",X"3B",X"11",X"10",X"8E",X"CD",X"66",X"C6",X"03",X"BD",X"38",
		X"50",X"BD",X"3B",X"24",X"8E",X"CD",X"3E",X"A6",X"C8",X"31",X"26",X"05",X"BF",X"BF",X"2A",X"20",
		X"03",X"BF",X"BF",X"2E",X"7E",X"43",X"3C",X"10",X"8E",X"CD",X"6C",X"20",X"36",X"34",X"12",X"10",
		X"8E",X"CF",X"AA",X"AE",X"C8",X"2D",X"8D",X"2B",X"25",X"0C",X"31",X"2E",X"10",X"8C",X"CF",X"F8",
		X"25",X"F4",X"1C",X"FE",X"35",X"92",X"31",X"3A",X"35",X"92",X"34",X"12",X"10",X"8E",X"CD",X"6C",
		X"AE",X"C8",X"2D",X"8D",X"0E",X"25",X"EF",X"31",X"2E",X"10",X"8C",X"CF",X"96",X"25",X"F4",X"1C",
		X"FE",X"35",X"92",X"34",X"36",X"1E",X"12",X"C6",X"04",X"8D",X"17",X"C1",X"04",X"26",X"02",X"84",
		X"0F",X"A1",X"A0",X"22",X"05",X"25",X"07",X"5A",X"26",X"EF",X"1C",X"FE",X"35",X"B6",X"1A",X"01",
		X"35",X"B6",X"8C",X"C0",X"00",X"25",X"04",X"BD",X"3C",X"7D",X"39",X"A6",X"80",X"39",X"8E",X"CC",
		X"16",X"BD",X"3C",X"8E",X"BD",X"3F",X"49",X"8E",X"26",X"43",X"20",X"02",X"C6",X"03",X"A7",X"25",
		X"E7",X"A4",X"AF",X"28",X"C6",X"02",X"E7",X"2E",X"C6",X"14",X"86",X"0A",X"30",X"2F",X"A7",X"80",
		X"5A",X"26",X"FB",X"8E",X"3F",X"75",X"AF",X"26",X"C6",X"0A",X"6F",X"21",X"E7",X"22",X"86",X"25",
		X"A7",X"23",X"AD",X"B8",X"06",X"25",X"15",X"10",X"AF",X"C8",X"36",X"ED",X"C8",X"32",X"86",X"03",
		X"BD",X"5D",X"9F",X"10",X"AE",X"C8",X"36",X"EC",X"C8",X"32",X"20",X"E6",X"6E",X"B8",X"0C",X"53",
		X"50",X"4C",X"41",X"54",X"2D",X"28",X"43",X"29",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",
		X"4C",X"49",X"41",X"4D",X"53",X"20",X"45",X"4C",X"45",X"43",X"54",X"52",X"4F",X"4E",X"49",X"43",
		X"53",X"20",X"49",X"4E",X"43",X"2E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"46",X"4A",X"7E",X"46",X"8B",X"7E",X"46",X"B0",X"7E",X"46",X"42",X"7E",X"46",X"84",X"7E",
		X"46",X"A9",X"7E",X"46",X"DB",X"7E",X"46",X"CE",X"46",X"FB",X"7E",X"46",X"D6",X"7E",X"46",X"C9",
		X"47",X"5F",X"34",X"67",X"10",X"8E",X"47",X"5F",X"20",X"06",X"34",X"67",X"10",X"8E",X"46",X"FB",
		X"1A",X"FF",X"F7",X"CA",X"01",X"8D",X"0E",X"35",X"E7",X"84",X"0F",X"81",X"0A",X"2F",X"02",X"86",
		X"0A",X"10",X"BE",X"BF",X"11",X"BF",X"CA",X"04",X"48",X"81",X"64",X"25",X"02",X"86",X"5A",X"10",
		X"AE",X"A6",X"EC",X"A1",X"FD",X"CA",X"06",X"10",X"BF",X"CA",X"02",X"C6",X"1A",X"F7",X"CA",X"00",
		X"5F",X"30",X"8B",X"39",X"34",X"67",X"CE",X"47",X"5F",X"20",X"05",X"34",X"67",X"CE",X"46",X"FB",
		X"1A",X"FF",X"FF",X"BF",X"11",X"F7",X"CA",X"01",X"CE",X"4E",X"71",X"33",X"C6",X"EE",X"C6",X"A6",
		X"C4",X"8D",X"BE",X"A6",X"C0",X"2A",X"F8",X"35",X"E7",X"34",X"67",X"CE",X"47",X"5F",X"20",X"05",
		X"34",X"67",X"CE",X"46",X"FB",X"1A",X"FF",X"FF",X"BF",X"11",X"F7",X"CA",X"01",X"44",X"44",X"44",
		X"44",X"8D",X"96",X"A6",X"61",X"8D",X"92",X"35",X"E7",X"7C",X"BF",X"36",X"20",X"03",X"7F",X"BF",
		X"36",X"CE",X"46",X"2C",X"20",X"0B",X"7C",X"BF",X"36",X"20",X"03",X"7F",X"BF",X"36",X"CE",X"46",
		X"23",X"10",X"8E",X"5C",X"9C",X"48",X"31",X"B6",X"AE",X"A1",X"EC",X"A1",X"7D",X"BF",X"36",X"27",
		X"01",X"5F",X"84",X"7F",X"AD",X"C4",X"6D",X"3E",X"2A",X"EE",X"39",X"47",X"C3",X"47",X"DA",X"47",
		X"F1",X"48",X"08",X"48",X"1F",X"48",X"36",X"48",X"4D",X"48",X"64",X"48",X"7B",X"48",X"92",X"48",
		X"A9",X"48",X"C0",X"48",X"D7",X"48",X"EE",X"49",X"05",X"49",X"1C",X"49",X"33",X"49",X"4A",X"49",
		X"61",X"49",X"78",X"49",X"88",X"49",X"9F",X"49",X"B6",X"49",X"CD",X"49",X"EB",X"4A",X"02",X"4A",
		X"19",X"4A",X"30",X"4A",X"47",X"4A",X"5E",X"4A",X"75",X"4A",X"8C",X"4A",X"A3",X"4A",X"BA",X"4A",
		X"D8",X"4A",X"EF",X"4B",X"06",X"4B",X"1D",X"4B",X"31",X"4B",X"3F",X"4B",X"56",X"4B",X"5F",X"4B",
		X"6F",X"4B",X"7F",X"4B",X"83",X"4B",X"93",X"4B",X"A3",X"4B",X"BA",X"4B",X"D1",X"4B",X"D7",X"4B",
		X"EE",X"4B",X"FA",X"4C",X"06",X"4C",X"12",X"4C",X"1E",X"4C",X"2A",X"4C",X"36",X"4C",X"42",X"4C",
		X"4E",X"4C",X"5A",X"4C",X"66",X"4C",X"6A",X"4C",X"76",X"4C",X"82",X"4C",X"8E",X"4C",X"9A",X"4C",
		X"A6",X"4C",X"B2",X"4C",X"BE",X"4C",X"CA",X"4C",X"D6",X"4C",X"E2",X"4C",X"EE",X"4C",X"FA",X"4D",
		X"0B",X"4B",X"EE",X"4D",X"17",X"4D",X"23",X"4D",X"2F",X"4C",X"2A",X"4D",X"3B",X"4D",X"47",X"4D",
		X"53",X"4D",X"7A",X"4D",X"8B",X"4D",X"97",X"4D",X"A3",X"4D",X"DA",X"4D",X"AF",X"4D",X"B7",X"4D",
		X"C3",X"4D",X"DA",X"4D",X"DA",X"4D",X"CA",X"4D",X"CE",X"4D",X"DA",X"4D",X"E6",X"4D",X"F7",X"4D",
		X"DA",X"4D",X"DA",X"03",X"07",X"11",X"11",X"10",X"10",X"01",X"10",X"10",X"01",X"10",X"10",X"01",
		X"10",X"10",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"03",X"07",X"00",X"11",X"10",X"01",
		X"11",X"10",X"11",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",
		X"10",X"03",X"07",X"11",X"11",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"11",X"00",X"01",
		X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"00",X"01",X"10",
		X"00",X"01",X"10",X"01",X"11",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"11",X"11",X"10",X"03",
		X"07",X"00",X"01",X"10",X"00",X"11",X"10",X"01",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",
		X"00",X"01",X"10",X"00",X"01",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"11",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"11",X"11",X"10",X"03",X"07",X"11",
		X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",
		X"10",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"00",X"01",X"10",X"00",X"11",X"00",X"01",
		X"10",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"03",X"07",X"11",X"11",X"10",
		X"11",X"00",X"10",X"11",X"00",X"10",X"01",X"11",X"00",X"11",X"00",X"10",X"11",X"00",X"10",X"11",
		X"11",X"00",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"11",X"10",
		X"00",X"00",X"10",X"00",X"00",X"10",X"11",X"11",X"10",X"03",X"07",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"07",X"11",X"11",X"10",X"11",X"11",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"10",X"01",
		X"10",X"10",X"01",X"10",X"10",X"01",X"10",X"03",X"07",X"11",X"11",X"00",X"11",X"01",X"10",X"11",
		X"01",X"10",X"11",X"11",X"00",X"11",X"01",X"10",X"11",X"01",X"10",X"11",X"11",X"00",X"03",X"07",
		X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",
		X"11",X"10",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"00",X"10",X"01",X"10",X"10",X"01",X"10",
		X"10",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"11",X"11",X"00",X"03",X"07",X"11",X"11",
		X"10",X"11",X"00",X"00",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"10",
		X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"11",X"00",X"11",X"00",
		X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",X"03",X"07",X"11",X"11",X"10",X"11",
		X"01",X"10",X"11",X"00",X"00",X"11",X"01",X"10",X"11",X"00",X"10",X"11",X"11",X"10",X"11",X"11",
		X"10",X"03",X"07",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"11",X"10",X"11",
		X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"02",X"07",X"11",X"00",X"11",X"00",X"11",X"00",
		X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"03",X"07",X"00",X"01",X"10",X"00",X"01",X"10",
		X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"10",X"01",X"10",X"11",X"11",X"10",X"03",
		X"07",X"11",X"00",X"10",X"11",X"01",X"00",X"11",X"10",X"00",X"11",X"10",X"00",X"11",X"11",X"00",
		X"11",X"01",X"10",X"11",X"00",X"10",X"03",X"07",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",
		X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"11",X"11",X"10",X"11",X"11",X"10",X"04",X"07",X"11",
		X"11",X"11",X"10",X"11",X"00",X"10",X"10",X"11",X"00",X"10",X"10",X"11",X"00",X"10",X"10",X"11",
		X"00",X"10",X"10",X"11",X"00",X"00",X"10",X"11",X"00",X"00",X"10",X"03",X"07",X"11",X"11",X"10",
		X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",
		X"00",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",
		X"11",X"00",X"10",X"11",X"11",X"10",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",
		X"10",X"11",X"11",X"10",X"11",X"11",X"10",X"11",X"00",X"00",X"11",X"00",X"00",X"11",X"00",X"00",
		X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"10",
		X"10",X"11",X"01",X"00",X"11",X"10",X"10",X"03",X"07",X"11",X"11",X"10",X"11",X"00",X"10",X"11",
		X"11",X"10",X"11",X"10",X"00",X"11",X"11",X"00",X"11",X"01",X"10",X"11",X"00",X"10",X"03",X"07",
		X"11",X"11",X"10",X"10",X"00",X"00",X"11",X"11",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"11",
		X"11",X"10",X"11",X"11",X"10",X"03",X"07",X"11",X"11",X"10",X"01",X"10",X"00",X"01",X"10",X"00",
		X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"01",X"10",X"00",X"03",X"07",X"11",X"00",
		X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"11",X"10",
		X"11",X"11",X"10",X"03",X"07",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",
		X"10",X"01",X"01",X"00",X"01",X"11",X"00",X"00",X"11",X"00",X"04",X"07",X"11",X"00",X"00",X"10",
		X"11",X"00",X"00",X"10",X"11",X"00",X"00",X"10",X"11",X"01",X"00",X"10",X"11",X"01",X"00",X"10",
		X"11",X"01",X"00",X"10",X"11",X"11",X"11",X"10",X"03",X"07",X"11",X"00",X"10",X"11",X"00",X"10",
		X"01",X"11",X"00",X"00",X"10",X"00",X"01",X"01",X"00",X"11",X"00",X"10",X"11",X"00",X"10",X"03",
		X"07",X"11",X"00",X"10",X"11",X"00",X"10",X"11",X"00",X"10",X"01",X"11",X"00",X"00",X"11",X"00",
		X"00",X"11",X"00",X"00",X"11",X"00",X"03",X"07",X"11",X"11",X"10",X"00",X"01",X"00",X"00",X"10",
		X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"11",X"11",X"10",X"11",X"11",X"10",X"03",X"06",X"00",
		X"00",X"00",X"00",X"10",X"00",X"01",X"10",X"00",X"11",X"11",X"10",X"01",X"10",X"00",X"00",X"10",
		X"00",X"03",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"03",
		X"07",X"01",X"11",X"00",X"10",X"00",X"10",X"10",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"07",X"10",X"10",X"10",X"10",X"10",X"00",X"10",X"02",
		X"07",X"00",X"10",X"01",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"01",X"00",X"00",X"10",X"02",
		X"07",X"10",X"00",X"01",X"00",X"00",X"10",X"00",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"01",
		X"02",X"10",X"10",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",
		X"00",X"01",X"00",X"02",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"11",X"00",X"03",X"07",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"01",X"00",X"00",X"10",
		X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"03",X"07",X"01",X"00",X"00",X"10",
		X"10",X"00",X"10",X"10",X"00",X"01",X"00",X"00",X"10",X"10",X"10",X"10",X"01",X"00",X"01",X"10",
		X"10",X"02",X"02",X"10",X"10",X"10",X"10",X"03",X"07",X"00",X"10",X"00",X"01",X"11",X"00",X"11",
		X"11",X"10",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"02",X"05",
		X"11",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"10",X"02",X"05",X"01",X"00",X"11",X"00",
		X"01",X"00",X"01",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"11",X"10",X"10",X"00",
		X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",X"10",X"02",X"05",
		X"10",X"10",X"10",X"10",X"11",X"10",X"00",X"10",X"00",X"10",X"02",X"05",X"11",X"10",X"10",X"00",
		X"11",X"10",X"00",X"10",X"11",X"10",X"02",X"05",X"11",X"10",X"10",X"00",X"11",X"10",X"10",X"10",
		X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"05",
		X"11",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"11",X"10",X"02",X"05",X"11",X"10",X"10",X"10",
		X"11",X"10",X"00",X"10",X"00",X"10",X"02",X"01",X"00",X"00",X"02",X"05",X"11",X"10",X"10",X"10",
		X"11",X"10",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",
		X"11",X"10",X"02",X"05",X"11",X"10",X"10",X"00",X"10",X"00",X"10",X"00",X"11",X"10",X"02",X"05",
		X"11",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"00",X"02",X"05",X"11",X"10",X"10",X"00",
		X"11",X"00",X"10",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"10",X"00",X"11",X"00",X"10",X"00",
		X"10",X"00",X"02",X"05",X"11",X"10",X"10",X"00",X"10",X"10",X"10",X"10",X"11",X"10",X"02",X"05",
		X"10",X"10",X"10",X"10",X"11",X"10",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"01",X"00",
		X"01",X"00",X"01",X"00",X"11",X"10",X"02",X"05",X"00",X"10",X"00",X"10",X"00",X"10",X"10",X"10",
		X"11",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"02",X"05",
		X"10",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"11",X"10",X"03",X"05",X"11",X"11",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"10",X"10",X"00",X"10",X"02",X"05",X"11",X"10",X"10",
		X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"10",X"10",X"11",X"10",X"10",
		X"00",X"10",X"00",X"02",X"05",X"11",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"00",X"10",X"02",
		X"05",X"11",X"10",X"10",X"10",X"11",X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"11",X"10",X"01",
		X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"02",X"05",X"10",X"10",X"10",X"10",X"10",X"10",X"10",
		X"10",X"11",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"10",X"10",X"01",X"00",X"01",X"00",X"53",
		X"50",X"4C",X"41",X"54",X"20",X"28",X"43",X"29",X"31",X"39",X"38",X"32",X"20",X"57",X"49",X"4C",
		X"4C",X"49",X"41",X"4D",X"53",X"20",X"49",X"4E",X"43",X"2E",X"03",X"05",X"10",X"00",X"10",X"10",
		X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"11",X"11",X"10",X"02",X"05",X"10",X"10",X"10",
		X"10",X"01",X"00",X"10",X"10",X"10",X"10",X"02",X"05",X"10",X"10",X"10",X"10",X"11",X"10",X"01",
		X"00",X"01",X"00",X"02",X"05",X"11",X"10",X"00",X"10",X"01",X"00",X"10",X"00",X"11",X"10",X"02",
		X"03",X"00",X"00",X"00",X"00",X"11",X"10",X"02",X"05",X"11",X"10",X"00",X"10",X"01",X"10",X"00",
		X"00",X"01",X"00",X"01",X"05",X"10",X"10",X"10",X"00",X"10",X"01",X"02",X"10",X"10",X"02",X"05",
		X"00",X"00",X"00",X"00",X"01",X"00",X"01",X"00",X"10",X"00",X"02",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"11",X"00",X"03",X"05",X"00",X"10",X"00",X"00",X"11",X"00",X"11",X"11",
		X"10",X"00",X"11",X"00",X"00",X"10",X"00",X"02",X"05",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"10",X"00",X"5A",X"07",X"5A",X"27",X"5A",X"46",X"5A",X"70",X"4F",X"EA",X"4F",X"D3",X"4F",
		X"BF",X"4F",X"9D",X"4F",X"89",X"4F",X"71",X"56",X"FE",X"56",X"F2",X"56",X"E9",X"56",X"C6",X"5B",
		X"43",X"5C",X"19",X"5B",X"F5",X"5B",X"DE",X"5B",X"BF",X"5B",X"23",X"5B",X"0A",X"5A",X"EB",X"58",
		X"D4",X"58",X"C6",X"58",X"B9",X"58",X"AC",X"58",X"A1",X"58",X"8B",X"58",X"6F",X"58",X"6A",X"5A",
		X"D5",X"5A",X"B2",X"5A",X"8A",X"58",X"66",X"58",X"62",X"58",X"5F",X"58",X"5C",X"58",X"59",X"58",
		X"56",X"58",X"41",X"58",X"31",X"58",X"18",X"58",X"02",X"57",X"F0",X"57",X"C2",X"57",X"B2",X"59",
		X"E4",X"59",X"C0",X"59",X"98",X"59",X"75",X"59",X"4C",X"59",X"27",X"59",X"08",X"58",X"EB",X"58",
		X"D9",X"4F",X"6D",X"57",X"DC",X"5B",X"A2",X"5B",X"81",X"5B",X"65",X"50",X"12",X"50",X"28",X"50",
		X"36",X"50",X"40",X"50",X"4A",X"50",X"55",X"50",X"65",X"50",X"7A",X"50",X"8E",X"50",X"90",X"50",
		X"97",X"50",X"A5",X"50",X"BC",X"50",X"D8",X"50",X"F0",X"50",X"FE",X"51",X"1A",X"51",X"25",X"51",
		X"2C",X"51",X"33",X"51",X"3D",X"51",X"4D",X"51",X"56",X"51",X"61",X"51",X"6C",X"51",X"7C",X"51",
		X"8C",X"51",X"95",X"51",X"9F",X"51",X"D6",X"51",X"E0",X"51",X"F2",X"52",X"01",X"52",X"12",X"52",
		X"22",X"52",X"2E",X"52",X"47",X"52",X"5C",X"52",X"6E",X"52",X"81",X"52",X"92",X"52",X"A6",X"52",
		X"BD",X"52",X"CD",X"52",X"E8",X"54",X"59",X"53",X"19",X"53",X"2A",X"53",X"3D",X"53",X"52",X"53",
		X"66",X"53",X"83",X"53",X"A6",X"53",X"C6",X"53",X"D8",X"53",X"F1",X"54",X"09",X"54",X"21",X"54",
		X"37",X"54",X"41",X"52",X"FF",X"54",X"69",X"54",X"87",X"54",X"AF",X"54",X"B2",X"54",X"BC",X"54",
		X"C2",X"54",X"DF",X"54",X"E7",X"55",X"00",X"55",X"22",X"55",X"3D",X"55",X"45",X"55",X"5B",X"55",
		X"67",X"55",X"7A",X"55",X"82",X"55",X"9F",X"56",X"7B",X"56",X"8E",X"56",X"B3",X"55",X"BD",X"55",
		X"DD",X"55",X"F0",X"56",X"08",X"56",X"18",X"56",X"4E",X"50",X"08",X"56",X"70",X"57",X"0E",X"57",
		X"16",X"57",X"1E",X"57",X"28",X"57",X"34",X"57",X"3E",X"57",X"49",X"57",X"56",X"57",X"63",X"57",
		X"74",X"00",X"00",X"5C",X"3A",X"56",X"D6",X"57",X"79",X"57",X"79",X"57",X"79",X"57",X"79",X"51",
		X"A6",X"51",X"AF",X"51",X"B9",X"51",X"C4",X"51",X"CC",X"57",X"7E",X"57",X"8F",X"00",X"76",X"5C",
		X"4E",X"5C",X"57",X"5C",X"59",X"5C",X"74",X"5C",X"7F",X"5C",X"89",X"5C",X"96",X"2C",X"00",X"00",
		X"80",X"12",X"0F",X"0B",X"0E",X"0A",X"2B",X"0F",X"17",X"0A",X"19",X"10",X"10",X"0A",X"0B",X"1E",
		X"0A",X"1E",X"12",X"0F",X"0A",X"1A",X"0B",X"1D",X"9D",X"0E",X"19",X"18",X"2B",X"1E",X"0A",X"16",
		X"19",X"1D",X"0F",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"12",X"0F",X"0B",X"8E",X"15",X"0F",X"0F",
		X"1A",X"0A",X"0B",X"0A",X"11",X"19",X"19",X"0E",X"0A",X"12",X"0F",X"0B",X"0E",X"0A",X"19",X"18",
		X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"1D",X"12",X"19",X"1F",X"16",X"0E",X"0F",X"1C",X"9D",X"1E",
		X"19",X"1F",X"11",X"12",X"0A",X"11",X"0F",X"1E",X"1E",X"13",X"18",X"11",X"0A",X"0B",X"12",X"0F",
		X"0B",X"0E",X"A7",X"16",X"19",X"19",X"15",X"2C",X"0A",X"0B",X"0A",X"0E",X"19",X"1F",X"0C",X"16",
		X"0F",X"1C",X"0A",X"12",X"0F",X"0B",X"0E",X"0F",X"1C",X"A8",X"23",X"19",X"1F",X"0A",X"18",X"0F",
		X"0F",X"0E",X"0A",X"0B",X"0A",X"12",X"0F",X"0B",X"0E",X"0A",X"1E",X"19",X"0A",X"1E",X"12",X"1C",
		X"19",X"21",X"0A",X"10",X"19",X"19",X"0E",X"A8",X"11",X"0B",X"17",X"0F",X"0A",X"19",X"20",X"0F",
		X"1C",X"8A",X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"0A",X"1E",X"0F",X"1D",X"1E",X"1D",X"0A",
		X"13",X"18",X"0E",X"13",X"0D",X"0B",X"1E",X"8F",X"0B",X"16",X"16",X"0A",X"1D",X"23",X"1D",X"1E",
		X"0F",X"17",X"1D",X"0A",X"11",X"99",X"1C",X"0B",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"8A",
		X"1C",X"19",X"17",X"0A",X"0F",X"1C",X"1C",X"19",X"1C",X"8A",X"0B",X"16",X"16",X"0A",X"1C",X"19",
		X"17",X"1D",X"0A",X"19",X"95",X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"1E",X"0A",X"10",X"19",
		X"16",X"16",X"19",X"21",X"9D",X"1A",X"1C",X"0F",X"1D",X"1D",X"0A",X"0B",X"0E",X"20",X"0B",X"18",
		X"0D",X"0F",X"0A",X"1E",X"19",X"0A",X"0F",X"22",X"13",X"9E",X"0A",X"1C",X"0B",X"17",X"0A",X"0F",
		X"1C",X"1C",X"19",X"1C",X"1D",X"0A",X"0E",X"0F",X"1E",X"0F",X"0D",X"1E",X"0F",X"8E",X"18",X"99",
		X"18",X"19",X"0A",X"0D",X"17",X"19",X"9D",X"0D",X"17",X"19",X"1D",X"0A",X"1C",X"0B",X"17",X"0A",
		X"0F",X"1C",X"1C",X"19",X"9C",X"10",X"1C",X"19",X"18",X"1E",X"0A",X"0E",X"19",X"19",X"1C",X"0A",
		X"17",X"1F",X"1D",X"1E",X"0A",X"0C",X"0F",X"0A",X"19",X"1A",X"0F",X"98",X"19",X"1C",X"0A",X"1E",
		X"0B",X"0C",X"16",X"0F",X"0A",X"1E",X"19",X"1A",X"0A",X"1C",X"0B",X"1D",X"13",X"0F",X"0E",X"0A",
		X"10",X"19",X"1C",X"0A",X"1E",X"0F",X"1D",X"9E",X"19",X"1C",X"0A",X"21",X"1C",X"13",X"1E",X"0F",
		X"0A",X"1A",X"1C",X"19",X"1E",X"0F",X"0D",X"1E",X"0A",X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",
		X"0D",X"19",X"16",X"19",X"1C",X"0A",X"1C",X"0B",X"17",X"0A",X"1E",X"0F",X"1D",X"9E",X"20",X"0F",
		X"1C",X"1E",X"13",X"0D",X"0B",X"16",X"0A",X"0C",X"0B",X"1C",X"1D",X"0A",X"13",X"18",X"0E",X"13",
		X"0D",X"0B",X"1E",X"0F",X"0A",X"0F",X"1C",X"1C",X"19",X"9C",X"1D",X"21",X"13",X"1E",X"0D",X"12",
		X"0A",X"1E",X"0F",X"1D",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"1F",X"9A",X"0B",X"0E",X"20",X"0B",
		X"18",X"0D",X"8F",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"0D",X"19",X"13",X"98",X"12",X"13",X"11",
		X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"16",X"0F",X"10",
		X"1E",X"0A",X"0D",X"19",X"13",X"98",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"0D",X"19",X"13",
		X"98",X"1D",X"16",X"0B",X"17",X"0A",X"1D",X"21",X"13",X"1E",X"0D",X"92",X"19",X"18",X"0F",X"0A",
		X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"1E",X"21",X"19",X"0A",
		X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"21",X"0B",X"16",X"15",
		X"0A",X"16",X"0F",X"10",X"9E",X"21",X"0B",X"16",X"15",X"0A",X"1C",X"13",X"11",X"12",X"9E",X"21",
		X"0B",X"16",X"15",X"0A",X"1F",X"9A",X"21",X"0B",X"16",X"15",X"0A",X"0E",X"19",X"21",X"98",X"1E",
		X"12",X"1C",X"19",X"21",X"0A",X"16",X"0F",X"10",X"9E",X"1E",X"12",X"1C",X"19",X"21",X"0A",X"1C",
		X"13",X"11",X"12",X"9E",X"1E",X"12",X"1C",X"19",X"21",X"0A",X"1F",X"9A",X"1E",X"12",X"1C",X"19",
		X"21",X"0A",X"0E",X"19",X"21",X"98",X"1D",X"19",X"1F",X"18",X"0E",X"0A",X"16",X"13",X"18",X"8F",
		X"0C",X"19",X"19",X"15",X"15",X"0F",X"0F",X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",
		X"16",X"9D",X"16",X"0F",X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",X"18",
		X"9D",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",
		X"18",X"9D",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"0D",X"19",X"13",
		X"18",X"9D",X"1A",X"0B",X"13",X"0E",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"9D",X"18",X"1F",
		X"17",X"0C",X"0F",X"1C",X"0A",X"19",X"10",X"0A",X"21",X"0B",X"20",X"0F",X"1D",X"0A",X"0D",X"19",
		X"17",X"1A",X"16",X"0F",X"1E",X"0F",X"8E",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"1E",X"13",X"17",
		X"0F",X"0A",X"13",X"18",X"0A",X"17",X"13",X"18",X"1F",X"1E",X"0F",X"9D",X"1E",X"19",X"1E",X"0B",
		X"16",X"0A",X"16",X"13",X"20",X"0F",X"1D",X"0A",X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"1E",X"19",
		X"1E",X"0B",X"16",X"0A",X"1D",X"13",X"18",X"11",X"16",X"0F",X"0A",X"1A",X"16",X"0B",X"23",X"0F",
		X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0E",X"1F",X"0B",X"16",X"0A",X"1A",X"16",X"0B",X"23",
		X"0F",X"9C",X"1E",X"19",X"1E",X"0B",X"16",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",X"1D",X"0A",
		X"1A",X"16",X"0B",X"23",X"0F",X"8E",X"0B",X"20",X"0F",X"1C",X"0B",X"11",X"0F",X"0A",X"1E",X"13",
		X"17",X"0F",X"0A",X"1A",X"0F",X"1C",X"0A",X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"11",X"0B",X"17",
		X"0F",X"0A",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",X"18",X"1E",X"9D",X"18",X"1F",X"17",
		X"0C",X"0F",X"1C",X"0A",X"19",X"10",X"0A",X"1D",X"0F",X"0D",X"19",X"18",X"0E",X"1D",X"0A",X"13",
		X"18",X"0A",X"0B",X"0A",X"21",X"0B",X"20",X"8F",X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"0A",
		X"18",X"1F",X"17",X"0C",X"0F",X"1C",X"0A",X"19",X"10",X"0A",X"16",X"13",X"20",X"0F",X"9D",X"12",
		X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"19",X"0A",X"0E",X"0B",X"1E",
		X"0F",X"0A",X"0B",X"16",X"16",X"19",X"21",X"0F",X"8E",X"1A",X"1C",X"13",X"0D",X"13",X"18",X"11",
		X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"13",X"19",X"98",X"0A",X"0A",X"0A",X"0A",X"16",X"0F",
		X"10",X"1E",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",
		X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"1D",X"16",X"19",X"1E",X"0A",X"1F",X"18",X"13",
		X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1D",X"16",X"19",X"1E",
		X"0A",X"1F",X"18",X"13",X"1E",X"9D",X"0A",X"0A",X"0A",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",
		X"1C",X"0F",X"1B",X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"0D",X"1C",X"0F",
		X"0E",X"13",X"9E",X"0A",X"0A",X"0A",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"1C",X"0F",X"1B",
		X"1F",X"13",X"1C",X"0F",X"0E",X"0A",X"10",X"19",X"1C",X"0A",X"0C",X"19",X"18",X"1F",X"1D",X"0A",
		X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0A",X"0A",X"0A",X"0A",X"17",X"13",X"18",X"13",X"17",X"1F",
		X"17",X"0A",X"1F",X"18",X"13",X"1E",X"1D",X"0A",X"10",X"19",X"1C",X"0A",X"0B",X"18",X"23",X"0A",
		X"0D",X"1C",X"0F",X"0E",X"13",X"9E",X"0E",X"13",X"10",X"10",X"13",X"0D",X"1F",X"16",X"1E",X"23",
		X"0A",X"19",X"10",X"0A",X"1A",X"16",X"0B",X"A3",X"16",X"0F",X"1E",X"1E",X"0F",X"1C",X"1D",X"0A",
		X"10",X"19",X"1C",X"0A",X"12",X"13",X"11",X"12",X"0F",X"1D",X"1E",X"0A",X"1D",X"0D",X"19",X"1C",
		X"8F",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"0A",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",
		X"0A",X"1D",X"0F",X"1E",X"1E",X"13",X"18",X"11",X"9D",X"0D",X"16",X"0F",X"0B",X"1C",X"0A",X"0C",
		X"19",X"19",X"15",X"15",X"0F",X"0F",X"1A",X"13",X"18",X"11",X"0A",X"1E",X"19",X"1E",X"0B",X"16",
		X"9D",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",X"1E",X"0B",X"0C",X"16",
		X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"0B",X"1F",X"1E",X"19",X"0A",X"0D",X"23",X"0D",X"16",
		X"8F",X"1D",X"0F",X"1E",X"0A",X"0B",X"1E",X"1E",X"1C",X"0B",X"0D",X"1E",X"0A",X"17",X"19",X"0E",
		X"0F",X"0A",X"17",X"0F",X"1D",X"1D",X"0B",X"11",X"8F",X"0F",X"22",X"1E",X"1C",X"0B",X"0A",X"16",
		X"13",X"10",X"0F",X"0A",X"0F",X"20",X"0F",X"1C",X"A3",X"1F",X"1D",X"0F",X"0A",X"2B",X"1A",X"16",
		X"0B",X"23",X"0F",X"1C",X"0A",X"01",X"0A",X"21",X"0B",X"16",X"15",X"2B",X"0A",X"1E",X"19",X"0A",
		X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"8A",X"1F",X"1D",X"0F",X"0A",X"2B",X"1A",X"16",X"0B",X"23",
		X"0F",X"1C",X"0A",X"01",X"0A",X"1E",X"12",X"1C",X"19",X"21",X"2B",X"0A",X"1E",X"19",X"0A",X"0D",
		X"12",X"0B",X"18",X"11",X"0F",X"0A",X"1E",X"12",X"0F",X"0A",X"20",X"0B",X"16",X"1F",X"8F",X"23",
		X"0F",X"9D",X"0B",X"0E",X"14",X"1F",X"1D",X"1E",X"17",X"0F",X"18",X"9E",X"16",X"0F",X"1E",X"1E",
		X"0F",X"9C",X"1F",X"1D",X"0F",X"0A",X"2B",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"01",X"0A",
		X"1E",X"12",X"1C",X"19",X"21",X"2B",X"0A",X"1E",X"19",X"0A",X"0F",X"18",X"1E",X"0F",X"9C",X"0A",
		X"10",X"0B",X"13",X"16",X"1F",X"1C",X"8F",X"10",X"0B",X"0D",X"1E",X"19",X"1C",X"23",X"0A",X"1D",
		X"0F",X"1E",X"1E",X"13",X"18",X"11",X"1D",X"0A",X"1C",X"0F",X"1D",X"1E",X"19",X"1C",X"0F",X"8E",
		X"0C",X"23",X"0A",X"19",X"1A",X"0F",X"18",X"13",X"18",X"11",X"0A",X"10",X"1C",X"19",X"18",X"1E",
		X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"19",X"1C",X"0A",X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1E",
		X"19",X"9A",X"0B",X"18",X"0E",X"0A",X"1E",X"1F",X"1C",X"18",X"13",X"18",X"11",X"0A",X"11",X"0B",
		X"17",X"0F",X"0A",X"19",X"18",X"0A",X"0B",X"18",X"0E",X"0A",X"19",X"10",X"90",X"0A",X"0D",X"16",
		X"0F",X"0B",X"1C",X"0F",X"8E",X"12",X"13",X"11",X"12",X"0A",X"1D",X"0D",X"19",X"1C",X"0F",X"0A",
		X"1E",X"0B",X"0C",X"16",X"0F",X"0A",X"1C",X"0F",X"1D",X"0F",X"9E",X"18",X"0F",X"1C",X"0E",X"0A",
		X"0C",X"0F",X"0B",X"1E",X"0F",X"1C",X"9D",X"1E",X"12",X"0F",X"0A",X"1D",X"1A",X"16",X"0B",X"1E",
		X"1E",X"13",X"18",X"11",X"0A",X"0F",X"16",X"13",X"1E",X"8F",X"0D",X"1C",X"0F",X"0E",X"13",X"1E",
		X"1D",X"8A",X"1F",X"1D",X"0F",X"0A",X"2B",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"01",X"0A",
		X"21",X"0B",X"16",X"15",X"2B",X"0A",X"1E",X"19",X"0A",X"0D",X"0F",X"18",X"1E",X"0F",X"9C",X"0F",
		X"18",X"1E",X"0F",X"1C",X"0A",X"16",X"13",X"18",X"0F",X"0A",X"0C",X"23",X"0A",X"1A",X"1C",X"0F",
		X"1D",X"1D",X"13",X"18",X"11",X"0A",X"0B",X"0E",X"20",X"0B",X"18",X"0D",X"8F",X"1A",X"1F",X"1E",
		X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"1D",X"0A",X"13",
		X"18",X"2D",X"2D",X"2D",X"0A",X"12",X"19",X"1E",X"0A",X"0E",X"19",X"11",X"8A",X"0F",X"18",X"1E",
		X"0F",X"1C",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"13",X"18",X"13",X"1E",X"13",X"0B",X"16",X"9D",
		X"23",X"19",X"1F",X"0A",X"0B",X"1C",X"0F",X"0A",X"18",X"19",X"21",X"0A",X"0B",X"0A",X"1D",X"1A",
		X"16",X"0B",X"1E",X"13",X"0B",X"1E",X"19",X"9C",X"17",X"0B",X"22",X"13",X"17",X"1F",X"17",X"0A",
		X"05",X"0A",X"0F",X"18",X"1E",X"1C",X"23",X"9D",X"1F",X"1D",X"0F",X"0A",X"26",X"21",X"0B",X"16",
		X"15",X"26",X"0A",X"1E",X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"0A",X"16",X"0F",X"1E",
		X"1E",X"0F",X"1C",X"0A",X"0A",X"0A",X"0A",X"26",X"1E",X"12",X"1C",X"19",X"21",X"26",X"0A",X"1E",
		X"19",X"0A",X"0F",X"18",X"1E",X"0F",X"1C",X"0A",X"16",X"0F",X"1E",X"1E",X"0F",X"9C",X"29",X"0D",
		X"2A",X"0A",X"01",X"09",X"08",X"02",X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",X"17",X"1D",X"0A",
		X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",X"0A",X"13",X"18",X"0D",X"AD",
		X"0A",X"0A",X"10",X"1C",X"0F",X"0F",X"0A",X"1A",X"16",X"0B",X"A3",X"1E",X"12",X"13",X"1D",X"0A",
		X"13",X"1D",X"0A",X"10",X"19",X"19",X"0E",X"0A",X"10",X"13",X"11",X"12",X"1E",X"AD",X"0E",X"0F",
		X"1D",X"13",X"11",X"18",X"0F",X"0E",X"0A",X"0C",X"23",X"0A",X"21",X"13",X"16",X"16",X"13",X"0B",
		X"17",X"1D",X"0A",X"0F",X"16",X"0F",X"0D",X"1E",X"1C",X"19",X"18",X"13",X"0D",X"1D",X"0A",X"13",
		X"18",X"0D",X"AD",X"0B",X"16",X"16",X"0A",X"1C",X"13",X"11",X"12",X"1E",X"1D",X"0A",X"1C",X"0F",
		X"1D",X"0F",X"1C",X"20",X"0F",X"8E",X"0D",X"1C",X"0F",X"0B",X"1E",X"1F",X"1C",X"0F",X"0A",X"10",
		X"0F",X"0B",X"1E",X"1F",X"1C",X"8F",X"0D",X"19",X"1C",X"18",X"0A",X"1D",X"1E",X"0B",X"16",X"15",
		X"0F",X"1C",X"0A",X"0B",X"1E",X"1E",X"0B",X"0D",X"95",X"18",X"0F",X"1C",X"0E",X"0A",X"12",X"1F",
		X"18",X"9E",X"13",X"18",X"1E",X"0F",X"1C",X"17",X"13",X"1D",X"1D",X"13",X"19",X"98",X"1E",X"1C",
		X"23",X"0A",X"1D",X"19",X"17",X"0F",X"0A",X"1A",X"19",X"1A",X"0D",X"19",X"1C",X"98",X"1A",X"16",
		X"0B",X"23",X"0F",X"1C",X"0A",X"81",X"1A",X"16",X"0B",X"23",X"0F",X"1C",X"0A",X"82",X"10",X"19",
		X"19",X"0E",X"0A",X"10",X"13",X"11",X"12",X"9E",X"0C",X"0B",X"18",X"0B",X"18",X"0B",X"0A",X"0C",
		X"1C",X"0B",X"21",X"96",X"1A",X"13",X"0F",X"0A",X"1A",X"1F",X"17",X"17",X"0F",X"96",X"10",X"13",
		X"1D",X"12",X"0A",X"10",X"13",X"0B",X"1D",X"0D",X"99",X"1E",X"19",X"17",X"0B",X"1E",X"19",X"0A",
		X"1E",X"1F",X"1D",X"1D",X"16",X"8F",X"0F",X"11",X"11",X"0A",X"0F",X"22",X"1A",X"16",X"19",X"1D",
		X"13",X"19",X"98",X"0C",X"0F",X"21",X"0B",X"1C",X"0F",X"0A",X"1E",X"12",X"0F",X"0A",X"12",X"13",
		X"1E",X"17",X"0B",X"98",X"1D",X"0D",X"19",X"1C",X"8F",X"21",X"0B",X"20",X"0F",X"8A",X"0D",X"12",
		X"19",X"19",X"1D",X"0F",X"0A",X"0D",X"12",X"0B",X"1C",X"0B",X"0D",X"1E",X"0F",X"1C",X"9D",X"17",
		X"19",X"20",X"0F",X"0A",X"21",X"0B",X"16",X"15",X"0A",X"14",X"19",X"23",X"1D",X"1E",X"13",X"0D",
		X"15",X"0A",X"1E",X"19",X"0A",X"1D",X"0F",X"16",X"0F",X"0D",X"1E",X"0A",X"1A",X"16",X"0B",X"23",
		X"0F",X"9C",X"1E",X"12",X"0F",X"0A",X"10",X"13",X"18",X"0F",X"1C",X"0A",X"1A",X"19",X"13",X"18",
		X"1E",X"9D",X"1D",X"1A",X"16",X"0B",X"1E",X"0A",X"21",X"13",X"1E",X"12",X"0A",X"1E",X"19",X"17",
		X"0B",X"1E",X"19",X"0F",X"1D",X"0A",X"26",X"0A",X"0F",X"11",X"11",X"9D",X"12",X"13",X"1E",X"0A",
		X"1E",X"12",X"0F",X"0A",X"0D",X"19",X"1C",X"18",X"0A",X"1D",X"1E",X"0B",X"16",X"15",X"0F",X"9C",
		X"1D",X"1A",X"16",X"0B",X"1E",X"0A",X"21",X"13",X"1E",X"12",X"0A",X"0C",X"0B",X"18",X"0B",X"18",
		X"0B",X"9D",X"1D",X"1A",X"16",X"0B",X"1E",X"0A",X"21",X"13",X"1E",X"12",X"0A",X"10",X"13",X"1D",
		X"12",X"0A",X"26",X"0A",X"15",X"0F",X"23",X"9D",X"1D",X"1A",X"16",X"0B",X"1E",X"0A",X"21",X"13",
		X"1E",X"12",X"0A",X"1A",X"13",X"0F",X"1D",X"0A",X"26",X"0A",X"1A",X"19",X"1A",X"0D",X"19",X"1C",
		X"98",X"1D",X"17",X"0B",X"0D",X"15",X"0A",X"0B",X"0A",X"18",X"0F",X"1C",X"0E",X"0A",X"10",X"19",
		X"9C",X"12",X"0B",X"17",X"17",X"0F",X"1C",X"0A",X"1E",X"12",X"0F",X"0A",X"12",X"13",X"1E",X"17",
		X"0B",X"18",X"0A",X"10",X"19",X"9C",X"02",X"05",X"80",X"04",X"00",X"80",X"05",X"00",X"80",X"07",
		X"05",X"80",X"01",X"05",X"00",X"80",X"01",X"00",X"00",X"80",X"02",X"00",X"00",X"00",X"A8",X"0F",
		X"22",X"1A",X"16",X"19",X"0E",X"0F",X"0A",X"1E",X"12",X"0F",X"0A",X"11",X"0B",X"1C",X"0C",X"0B",
		X"11",X"0F",X"0A",X"0D",X"1C",X"0F",X"0B",X"1E",X"1F",X"1C",X"8F",X"1D",X"1A",X"16",X"0B",X"1E",
		X"0A",X"1E",X"12",X"0F",X"0A",X"19",X"1E",X"12",X"0F",X"1C",X"0A",X"1A",X"16",X"0B",X"23",X"0F",
		X"9C",X"12",X"0F",X"0B",X"0E",X"0A",X"12",X"19",X"18",X"0D",X"12",X"99",X"1E",X"0B",X"18",X"23",
		X"0B",X"0A",X"1E",X"19",X"19",X"1E",X"1D",X"13",X"8F",X"17",X"0B",X"1C",X"0D",X"0A",X"1E",X"12",
		X"0F",X"0A",X"1D",X"16",X"19",X"8C",X"12",X"0B",X"1C",X"1C",X"23",X"0A",X"1E",X"12",X"0F",X"0A",
		X"12",X"19",X"19",X"8E",X"16",X"13",X"20",X"0F",X"9D",X"1E",X"12",X"0F",X"0A",X"1C",X"1F",X"16",
		X"0F",X"1D",X"0A",X"19",X"10",X"0A",X"1D",X"1A",X"16",X"0B",X"9E",X"23",X"19",X"1F",X"0A",X"0B",
		X"1C",X"0F",X"0A",X"19",X"18",X"0F",X"0A",X"19",X"10",X"0A",X"1D",X"1A",X"16",X"0B",X"1E",X"2B",
		X"1D",X"0A",X"0F",X"16",X"13",X"1E",X"0F",X"AF",X"23",X"19",X"1F",X"0A",X"10",X"13",X"11",X"12",
		X"1E",X"0A",X"1E",X"19",X"0A",X"21",X"13",X"18",X"2C",X"0A",X"0B",X"20",X"19",X"13",X"0E",X"0A",
		X"0E",X"0F",X"10",X"0F",X"0B",X"1E",X"AD",X"11",X"19",X"0A",X"11",X"1C",X"0B",X"0C",X"0A",X"1D",
		X"19",X"17",X"0F",X"0A",X"10",X"19",X"19",X"0E",X"0A",X"1E",X"12",X"0B",X"1E",X"0A",X"10",X"0B",
		X"16",X"16",X"1D",X"0A",X"13",X"18",X"0A",X"1C",X"19",X"21",X"1D",X"AF",X"1E",X"12",X"0F",X"18",
		X"0A",X"1E",X"12",X"1C",X"19",X"21",X"0A",X"13",X"1E",X"0A",X"1B",X"1F",X"13",X"0D",X"15",X"2C",
		X"0A",X"0B",X"18",X"0E",X"0A",X"1D",X"1A",X"16",X"0B",X"1E",X"0A",X"23",X"19",X"1F",X"1C",X"0A",
		X"10",X"19",X"0F",X"1D",X"AD",X"13",X"10",X"0A",X"12",X"13",X"1E",X"0A",X"0C",X"23",X"0A",X"10",
		X"19",X"19",X"0E",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"12",X"0F",X"0B",X"0E",X"0A",X"21",X"13",
		X"16",X"16",X"0A",X"1C",X"19",X"16",X"16",X"AF",X"23",X"19",X"1F",X"2B",X"1C",X"0F",X"0A",X"12",
		X"0F",X"16",X"1A",X"16",X"0F",X"1D",X"1D",X"0A",X"1E",X"12",X"0F",X"18",X"0A",X"1F",X"18",X"1E",
		X"13",X"16",X"0A",X"23",X"19",X"1F",X"2B",X"1C",X"0F",X"0A",X"21",X"12",X"19",X"16",X"0F",X"AD",
		X"11",X"19",X"0A",X"1D",X"1A",X"16",X"0B",X"1E",X"1E",X"0F",X"1C",X"0A",X"18",X"0F",X"1C",X"0E",
		X"1D",X"0A",X"10",X"19",X"1C",X"0A",X"12",X"13",X"11",X"12",X"0F",X"1C",X"0A",X"1D",X"0D",X"19",
		X"1C",X"0F",X"1D",X"AF",X"1A",X"13",X"0D",X"15",X"0A",X"1F",X"1A",X"0A",X"10",X"19",X"19",X"0E",
		X"0A",X"10",X"16",X"23",X"13",X"18",X"11",X"0A",X"10",X"1C",X"19",X"17",X"0A",X"1E",X"12",X"0F",
		X"0A",X"0E",X"19",X"19",X"1C",X"1D",X"AD",X"19",X"18",X"0A",X"0F",X"18",X"1E",X"0F",X"1C",X"13",
		X"18",X"11",X"2C",X"0A",X"1E",X"12",X"0F",X"0A",X"0E",X"19",X"19",X"1C",X"0A",X"23",X"19",X"1F",
		X"0A",X"0D",X"12",X"19",X"19",X"1D",X"8F",X"21",X"13",X"16",X"16",X"0A",X"10",X"16",X"0B",X"1D",
		X"12",X"0A",X"0C",X"1C",X"13",X"11",X"12",X"1E",X"0A",X"1C",X"0F",X"0E",X"0A",X"0B",X"18",X"0E",
		X"0A",X"11",X"16",X"19",X"21",X"AF",X"23",X"19",X"1F",X"0A",X"0D",X"12",X"0B",X"18",X"11",X"0F",
		X"0A",X"13",X"1E",X"0A",X"21",X"13",X"1E",X"12",X"0A",X"1E",X"12",X"0F",X"0A",X"1D",X"1E",X"13",
		X"0D",X"15",X"0A",X"17",X"0B",X"1C",X"15",X"0F",X"0E",X"0A",X"2B",X"17",X"19",X"20",X"0F",X"AB",
		X"0B",X"18",X"0E",X"0A",X"0D",X"19",X"17",X"0F",X"0A",X"19",X"1F",X"1E",X"0A",X"1F",X"1D",X"13",
		X"18",X"11",X"0A",X"2B",X"1E",X"12",X"1C",X"19",X"21",X"AB",X"1A",X"0B",X"1D",X"1D",X"0A",X"1E",
		X"12",X"1C",X"19",X"1F",X"11",X"12",X"0A",X"1E",X"12",X"0F",X"0A",X"0E",X"19",X"19",X"1C",X"1D",
		X"0A",X"0C",X"23",X"0A",X"0D",X"0B",X"1E",X"0D",X"12",X"13",X"18",X"11",X"0A",X"15",X"0F",X"23",
		X"1D",X"AF",X"0B",X"18",X"0E",X"0A",X"1C",X"0F",X"0B",X"0D",X"12",X"0A",X"1E",X"12",X"0F",X"0A",
		X"19",X"1E",X"12",X"0F",X"1C",X"0A",X"1D",X"13",X"0E",X"0F",X"0A",X"21",X"13",X"1E",X"12",X"0A",
		X"0F",X"0B",X"1D",X"0F",X"AD",X"23",X"19",X"1F",X"1C",X"0A",X"0F",X"18",X"0F",X"17",X"13",X"0F",
		X"1D",X"0A",X"0B",X"1C",X"0F",X"0A",X"18",X"0B",X"1D",X"1E",X"A3",X"1E",X"12",X"0F",X"23",X"0A",
		X"21",X"13",X"16",X"16",X"0A",X"0D",X"12",X"0B",X"1D",X"0F",X"0A",X"0B",X"18",X"0E",X"0A",X"0C",
		X"19",X"1E",X"12",X"0F",X"1C",X"0A",X"23",X"19",X"1F",X"AF",X"0C",X"0F",X"21",X"0B",X"1C",X"0F",
		X"0A",X"19",X"10",X"0A",X"1D",X"1A",X"0F",X"0F",X"0E",X"23",X"0A",X"12",X"13",X"1E",X"0A",X"17",
		X"0F",X"18",X"AC",X"1A",X"0F",X"0F",X"16",X"1D",X"2C",X"0A",X"0B",X"18",X"0E",X"0A",X"1A",X"19",
		X"1A",X"0D",X"19",X"1C",X"18",X"0A",X"1D",X"1E",X"0B",X"16",X"15",X"0F",X"1C",X"1D",X"0A",X"1E",
		X"19",X"19",X"AD",X"1E",X"12",X"0F",X"0A",X"11",X"0B",X"1C",X"0C",X"0B",X"11",X"0F",X"0A",X"0D",
		X"1C",X"0F",X"0B",X"1E",X"1F",X"1C",X"0F",X"1D",X"0A",X"12",X"19",X"1A",X"0A",X"0B",X"18",X"0E",
		X"0A",X"14",X"1F",X"17",X"9A",X"0E",X"19",X"18",X"2B",X"1E",X"0A",X"16",X"0F",X"1E",X"0A",X"1E",
		X"12",X"0F",X"17",X"0A",X"11",X"0F",X"1E",X"0A",X"1E",X"19",X"19",X"0A",X"18",X"0F",X"0B",X"1C",
		X"AC",X"19",X"18",X"0F",X"0A",X"12",X"13",X"1E",X"0A",X"21",X"13",X"16",X"16",X"0A",X"1D",X"16",
		X"19",X"21",X"0A",X"1E",X"12",X"0F",X"17",X"0A",X"0E",X"19",X"21",X"18",X"0A",X"0B",X"0A",X"0C",
		X"13",X"9E",X"1E",X"21",X"19",X"0A",X"12",X"13",X"1E",X"1D",X"0A",X"23",X"19",X"1F",X"2B",X"1C",
		X"0F",X"0A",X"13",X"18",X"0A",X"1E",X"12",X"0F",X"0A",X"0D",X"16",X"0F",X"0B",X"1C",X"AD",X"23",
		X"19",X"1F",X"1C",X"0A",X"10",X"0F",X"16",X"16",X"19",X"21",X"0A",X"1A",X"16",X"0B",X"23",X"0F",
		X"1C",X"0A",X"0B",X"1E",X"0A",X"23",X"19",X"1F",X"1C",X"0A",X"1D",X"13",X"0E",X"8F",X"0D",X"0B",
		X"18",X"0A",X"0B",X"13",X"0E",X"0A",X"23",X"19",X"1F",X"2C",X"0A",X"19",X"1C",X"0A",X"0C",X"0F",
		X"1E",X"1C",X"0B",X"23",X"AF",X"13",X"1E",X"2B",X"1D",X"0A",X"1C",X"19",X"1F",X"11",X"12",X"0A",
		X"21",X"12",X"0F",X"18",X"0A",X"23",X"19",X"1F",X"2B",X"1C",X"0F",X"0A",X"18",X"19",X"1E",X"0A",
		X"10",X"1C",X"13",X"0F",X"18",X"0E",X"16",X"23",X"AC",X"0C",X"1F",X"1E",X"0A",X"23",X"19",X"1F",
		X"0A",X"11",X"0F",X"1E",X"0A",X"17",X"19",X"1C",X"0F",X"0A",X"1A",X"19",X"13",X"18",X"1E",X"1D",
		X"0A",X"1E",X"12",X"0B",X"1E",X"0A",X"21",X"0B",X"23",X"AD",X"02",X"0A",X"12",X"13",X"1E",X"1D",
		X"0A",X"15",X"13",X"16",X"16",X"0A",X"0D",X"1C",X"0F",X"0B",X"1E",X"1F",X"1C",X"8F",X"0A",X"1E",
		X"19",X"0A",X"1D",X"1E",X"0B",X"1C",X"9E",X"19",X"9C",X"13",X"18",X"1D",X"0F",X"1C",X"1E",X"0A",
		X"0B",X"0E",X"0E",X"13",X"1E",X"13",X"19",X"18",X"0B",X"16",X"0A",X"0D",X"19",X"13",X"18",X"1D",
		X"0A",X"10",X"19",X"9C",X"30",X"0E",X"1F",X"0B",X"16",X"0A",X"1A",X"16",X"0B",X"23",X"B0",X"1C",
		X"0F",X"0B",X"0E",X"23",X"0A",X"10",X"19",X"1C",X"8A",X"30",X"1D",X"13",X"18",X"11",X"16",X"0F",
		X"0A",X"1A",X"16",X"0B",X"23",X"B0",X"1A",X"1C",X"0F",X"1D",X"1D",X"8A",X"5C",X"C4",X"5C",X"D0",
		X"5C",X"D8",X"5C",X"E0",X"5C",X"E4",X"5C",X"F4",X"5C",X"FC",X"5D",X"00",X"5D",X"04",X"5D",X"08",
		X"5D",X"18",X"5D",X"28",X"5D",X"3C",X"5D",X"40",X"5D",X"48",X"5D",X"4C",X"5D",X"4C",X"5D",X"54",
		X"5D",X"64",X"5D",X"7C",X"3E",X"50",X"09",X"99",X"36",X"90",X"0A",X"33",X"2E",X"A0",X"8B",X"33",
		X"2A",X"80",X"0D",X"99",X"30",X"80",X"8C",X"99",X"21",X"80",X"0E",X"99",X"37",X"80",X"8C",X"99",
		X"36",X"80",X"8F",X"22",X"36",X"80",X"0F",X"22",X"28",X"90",X"12",X"22",X"17",X"A0",X"10",X"99",
		X"17",X"A8",X"91",X"99",X"3A",X"80",X"13",X"33",X"24",X"B0",X"94",X"33",X"3A",X"20",X"95",X"88",
		X"2F",X"10",X"A3",X"99",X"2F",X"10",X"AF",X"99",X"23",X"D7",X"42",X"BB",X"5E",X"D7",X"45",X"BB",
		X"25",X"DF",X"43",X"44",X"34",X"E7",X"8B",X"11",X"28",X"16",X"40",X"BB",X"16",X"C0",X"42",X"33",
		X"6D",X"C0",X"46",X"33",X"20",X"D0",X"C7",X"33",X"30",X"80",X"45",X"22",X"4F",X"80",X"48",X"22",
		X"27",X"A0",X"3C",X"22",X"19",X"B0",X"4A",X"22",X"23",X"C0",X"CB",X"22",X"21",X"80",X"C9",X"99",
		X"24",X"60",X"23",X"33",X"59",X"60",X"CC",X"33",X"2A",X"40",X"CD",X"88",X"3A",X"2A",X"4E",X"11",
		X"31",X"60",X"CF",X"22",X"10",X"30",X"53",X"11",X"10",X"40",X"54",X"11",X"10",X"50",X"5B",X"11",
		X"10",X"60",X"D5",X"11",X"24",X"57",X"7D",X"11",X"36",X"57",X"7C",X"55",X"5A",X"57",X"77",X"11",
		X"49",X"77",X"78",X"11",X"26",X"97",X"79",X"11",X"3D",X"A7",X"FA",X"77",X"2E",X"77",X"7B",X"11",
		X"4D",X"77",X"FA",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7E",X"E6",X"AA",X"7E",X"7F",X"1D",X"7E",X"E3",X"40",X"7E",X"D6",X"76",X"7E",X"D6",X"C5",X"7E",
		X"D6",X"BA",X"7E",X"D6",X"F6",X"E6",X"96",X"7E",X"79",X"75",X"7E",X"6E",X"C3",X"7E",X"84",X"4A",
		X"7E",X"6C",X"01",X"7E",X"6D",X"26",X"7E",X"74",X"AF",X"7E",X"6B",X"F3",X"7E",X"8D",X"DD",X"34",
		X"04",X"DC",X"1F",X"53",X"C5",X"09",X"26",X"05",X"53",X"46",X"56",X"20",X"09",X"53",X"C5",X"09",
		X"26",X"02",X"27",X"F5",X"44",X"56",X"DD",X"1F",X"35",X"84",X"39",X"2A",X"FD",X"E6",X"15",X"C1",
		X"F0",X"27",X"F7",X"6C",X"02",X"1F",X"89",X"EB",X"15",X"34",X"07",X"1A",X"F0",X"E7",X"15",X"CC",
		X"AA",X"CC",X"FD",X"CA",X"04",X"10",X"AE",X"1A",X"EC",X"3E",X"FD",X"CA",X"06",X"10",X"BF",X"CA",
		X"02",X"C6",X"02",X"F7",X"CA",X"00",X"E6",X"61",X"2A",X"34",X"A6",X"62",X"80",X"06",X"2B",X"01",
		X"4F",X"AB",X"3E",X"27",X"02",X"2A",X"05",X"86",X"F0",X"A7",X"15",X"4F",X"B7",X"CA",X"06",X"E6",
		X"3E",X"EB",X"62",X"34",X"04",X"A0",X"3E",X"40",X"8B",X"AA",X"C6",X"CC",X"FD",X"CA",X"02",X"A6",
		X"63",X"81",X"06",X"2A",X"02",X"86",X"06",X"E6",X"17",X"FD",X"CA",X"04",X"20",X"26",X"86",X"90",
		X"A0",X"62",X"27",X"02",X"2A",X"05",X"86",X"F0",X"A7",X"15",X"4F",X"A1",X"3E",X"23",X"02",X"A6",
		X"3E",X"B7",X"CA",X"06",X"CC",X"AA",X"CC",X"FD",X"CA",X"02",X"A6",X"62",X"E6",X"17",X"FD",X"CA",
		X"04",X"4A",X"34",X"02",X"E6",X"15",X"C1",X"F0",X"27",X"05",X"C6",X"07",X"F7",X"CA",X"00",X"86",
		X"01",X"35",X"04",X"B7",X"CA",X"06",X"F7",X"CA",X"04",X"7F",X"CA",X"01",X"C6",X"12",X"F7",X"CA",
		X"00",X"35",X"87",X"AE",X"49",X"BD",X"D7",X"84",X"BD",X"DC",X"73",X"10",X"AE",X"47",X"10",X"AE",
		X"35",X"10",X"AF",X"47",X"20",X"1D",X"8E",X"E6",X"7E",X"BD",X"E6",X"AA",X"86",X"08",X"20",X"02",
		X"86",X"0A",X"AE",X"49",X"E6",X"03",X"BD",X"D7",X"84",X"BD",X"DC",X"73",X"10",X"AE",X"47",X"C5",
		X"03",X"26",X"07",X"BD",X"5D",X"BF",X"C6",X"04",X"3D",X"48",X"E6",X"39",X"C1",X"40",X"27",X"02",
		X"6C",X"2C",X"BD",X"5F",X"31",X"97",X"3C",X"BD",X"5D",X"BF",X"8A",X"3F",X"A7",X"1D",X"BD",X"5D",
		X"BF",X"4F",X"D6",X"1F",X"CA",X"0F",X"2A",X"02",X"4A",X"53",X"ED",X"1E",X"A6",X"35",X"81",X"4D",
		X"24",X"04",X"6A",X"1C",X"60",X"1D",X"5F",X"ED",X"11",X"ED",X"15",X"A6",X"37",X"A7",X"13",X"ED",
		X"17",X"10",X"8E",X"5F",X"52",X"96",X"3C",X"31",X"A6",X"10",X"AF",X"08",X"BD",X"D8",X"C6",X"A6",
		X"15",X"81",X"06",X"25",X"06",X"AB",X"B4",X"81",X"90",X"23",X"02",X"6F",X"11",X"9F",X"2E",X"AF",
		X"4B",X"86",X"14",X"BD",X"D6",X"BA",X"AE",X"47",X"A6",X"19",X"81",X"40",X"27",X"02",X"6F",X"0C",
		X"86",X"0F",X"BD",X"D6",X"BA",X"AE",X"4B",X"A6",X"11",X"26",X"F5",X"BD",X"D7",X"7D",X"7E",X"D6",
		X"C5",X"34",X"06",X"9E",X"30",X"26",X"01",X"3F",X"EC",X"84",X"DD",X"30",X"DC",X"2E",X"ED",X"84",
		X"4F",X"5F",X"A7",X"02",X"ED",X"1C",X"ED",X"1E",X"A7",X"04",X"A7",X"05",X"A7",X"0C",X"EF",X"0A",
		X"35",X"86",X"1C",X"C8",X"1D",X"D6",X"1D",X"12",X"1D",X"74",X"1E",X"1E",X"1E",X"58",X"C3",X"D6",
		X"D7",X"E8",X"D9",X"C9",X"C7",X"C8",X"E3",X"40",X"4D",X"C3",X"5D",X"40",X"F1",X"F9",X"F8",X"F2",
		X"40",X"E6",X"C9",X"D3",X"D3",X"C9",X"C1",X"D4",X"E2",X"40",X"C5",X"D3",X"C5",X"C3",X"E3",X"D9",
		X"D6",X"D5",X"C9",X"C3",X"E2",X"6B",X"40",X"C9",X"D5",X"C3",X"4B",X"00",X"39",X"6F",X"48",X"6F",
		X"47",X"86",X"05",X"BD",X"D6",X"BA",X"B6",X"99",X"84",X"BB",X"99",X"CC",X"27",X"29",X"2B",X"10",
		X"A6",X"48",X"27",X"ED",X"6A",X"48",X"26",X"E9",X"A6",X"49",X"C6",X"FF",X"8D",X"2B",X"20",X"E1",
		X"A6",X"48",X"26",X"DD",X"6A",X"47",X"2A",X"04",X"86",X"03",X"A7",X"47",X"A6",X"47",X"C6",X"14",
		X"E7",X"48",X"5F",X"A7",X"49",X"20",X"E5",X"A6",X"48",X"27",X"0A",X"A6",X"49",X"81",X"04",X"27",
		X"CF",X"C6",X"FF",X"8D",X"04",X"86",X"04",X"20",X"E5",X"8E",X"5F",X"EC",X"48",X"48",X"30",X"86",
		X"A6",X"84",X"5D",X"26",X"02",X"E6",X"03",X"AE",X"01",X"7E",X"46",X"2C",X"D2",X"31",X"EC",X"22",
		X"D1",X"37",X"EC",X"22",X"D0",X"26",X"EC",X"22",X"CF",X"35",X"EC",X"22",X"CE",X"33",X"EC",X"11",
		X"BD",X"5F",X"31",X"CC",X"32",X"15",X"ED",X"08",X"6F",X"11",X"9F",X"2E",X"AF",X"47",X"AE",X"47",
		X"A6",X"11",X"27",X"22",X"6F",X"D8",X"0D",X"BD",X"5D",X"AD",X"26",X"2B",X"DE",X"1C",X"AE",X"47",
		X"96",X"CB",X"27",X"0C",X"A6",X"05",X"81",X"02",X"27",X"15",X"6A",X"4C",X"26",X"11",X"20",X"17",
		X"6A",X"4B",X"27",X"5A",X"20",X"09",X"A6",X"D8",X"0D",X"26",X"21",X"96",X"CB",X"26",X"1D",X"86",
		X"04",X"8E",X"60",X"0E",X"7E",X"D6",X"BC",X"DE",X"1C",X"AE",X"47",X"A6",X"04",X"4C",X"8D",X"4F",
		X"86",X"64",X"A7",X"4B",X"A6",X"05",X"81",X"03",X"27",X"1E",X"20",X"E3",X"AE",X"47",X"5F",X"A6",
		X"4A",X"BB",X"32",X"19",X"A7",X"13",X"ED",X"17",X"BD",X"D8",X"C6",X"A6",X"49",X"BB",X"32",X"17",
		X"ED",X"15",X"ED",X"11",X"8D",X"44",X"20",X"D8",X"86",X"08",X"BD",X"D6",X"BA",X"86",X"04",X"AE",
		X"47",X"8D",X"1C",X"86",X"08",X"BD",X"D6",X"BA",X"86",X"02",X"AE",X"47",X"20",X"C0",X"86",X"64",
		X"A7",X"4B",X"A6",X"04",X"4A",X"2A",X"04",X"6F",X"15",X"20",X"A4",X"8D",X"02",X"20",X"B1",X"1A",
		X"50",X"A7",X"05",X"C6",X"05",X"3D",X"10",X"8E",X"32",X"15",X"31",X"A5",X"A6",X"49",X"AB",X"22",
		X"A7",X"15",X"A6",X"4A",X"AB",X"24",X"A7",X"17",X"1C",X"AF",X"86",X"0A",X"A7",X"4C",X"39",X"1D",
		X"D0",X"50",X"1D",X"E7",X"6D",X"D0",X"50",X"6D",X"E7",X"43",X"3D",X"5A",X"00",X"00",X"BD",X"5D",
		X"BF",X"C6",X"03",X"3D",X"C6",X"05",X"3D",X"10",X"8E",X"60",X"BF",X"31",X"A5",X"EC",X"A4",X"DD",
		X"BD",X"BE",X"99",X"86",X"A6",X"11",X"27",X"07",X"BD",X"89",X"35",X"A1",X"22",X"25",X"0E",X"BE",
		X"99",X"CE",X"A6",X"11",X"27",X"15",X"BD",X"89",X"35",X"A1",X"22",X"24",X"0E",X"31",X"25",X"10",
		X"8C",X"60",X"CD",X"25",X"D8",X"10",X"8E",X"60",X"BF",X"20",X"D2",X"EC",X"23",X"26",X"20",X"86",
		X"04",X"BD",X"E9",X"72",X"86",X"05",X"BD",X"D6",X"BA",X"EC",X"9F",X"34",X"0E",X"A7",X"C8",X"35",
		X"E7",X"C8",X"37",X"CC",X"61",X"61",X"ED",X"C8",X"38",X"CC",X"34",X"D3",X"7E",X"85",X"A6",X"ED",
		X"47",X"6F",X"49",X"E6",X"49",X"5C",X"BE",X"34",X"0E",X"E1",X"01",X"22",X"29",X"E7",X"49",X"6A",
		X"48",X"A6",X"84",X"1A",X"50",X"30",X"02",X"BF",X"CA",X"02",X"FD",X"CA",X"06",X"EC",X"47",X"FD",
		X"CA",X"04",X"86",X"02",X"B7",X"CA",X"00",X"1C",X"AF",X"86",X"02",X"8E",X"61",X"33",X"7E",X"D6",
		X"BC",X"CC",X"44",X"37",X"ED",X"47",X"BD",X"D7",X"3C",X"34",X"0E",X"94",X"96",X"77",X"2B",X"04",
		X"9F",X"77",X"20",X"02",X"9F",X"79",X"86",X"0E",X"A7",X"19",X"A6",X"47",X"5F",X"ED",X"11",X"ED",
		X"15",X"A6",X"48",X"ED",X"17",X"81",X"37",X"26",X"02",X"80",X"02",X"A7",X"13",X"E7",X"C8",X"1E",
		X"E7",X"C8",X"19",X"E7",X"4C",X"BD",X"D8",X"C6",X"AF",X"47",X"9F",X"2A",X"DC",X"EB",X"ED",X"4D",
		X"ED",X"C8",X"11",X"DC",X"EE",X"ED",X"4F",X"ED",X"C8",X"13",X"BD",X"63",X"4B",X"0C",X"B7",X"96",
		X"B7",X"44",X"24",X"0B",X"DC",X"EB",X"E3",X"4D",X"ED",X"4D",X"ED",X"C8",X"11",X"20",X"09",X"DC",
		X"EE",X"E3",X"4F",X"ED",X"4F",X"ED",X"C8",X"13",X"BE",X"99",X"86",X"BD",X"5D",X"BF",X"2B",X"03",
		X"BE",X"99",X"CE",X"AF",X"4A",X"86",X"02",X"A7",X"C8",X"1A",X"AE",X"47",X"E6",X"C8",X"1E",X"E1",
		X"C8",X"19",X"26",X"2B",X"6A",X"C8",X"21",X"26",X"0A",X"EC",X"C8",X"13",X"ED",X"4F",X"EC",X"C8",
		X"11",X"ED",X"4D",X"10",X"AE",X"06",X"10",X"2A",X"01",X"DA",X"6F",X"06",X"AE",X"2A",X"8C",X"99",
		X"91",X"10",X"27",X"01",X"50",X"8C",X"99",X"D9",X"10",X"27",X"01",X"49",X"7E",X"63",X"D4",X"E7",
		X"C8",X"19",X"6F",X"06",X"BE",X"99",X"86",X"E6",X"49",X"C5",X"02",X"26",X"07",X"C5",X"01",X"27",
		X"05",X"BE",X"99",X"CE",X"AF",X"4A",X"8E",X"E6",X"81",X"BD",X"E6",X"AA",X"EC",X"4F",X"47",X"56",
		X"47",X"56",X"DD",X"43",X"47",X"56",X"E3",X"4F",X"ED",X"C8",X"13",X"DC",X"43",X"E3",X"4F",X"43",
		X"50",X"82",X"FF",X"ED",X"4F",X"EC",X"4D",X"47",X"56",X"47",X"56",X"DD",X"43",X"47",X"56",X"E3",
		X"4D",X"ED",X"C8",X"11",X"DC",X"43",X"E3",X"4D",X"43",X"50",X"82",X"FF",X"ED",X"4D",X"C6",X"03",
		X"E7",X"C8",X"1D",X"20",X"03",X"BD",X"63",X"4B",X"86",X"0A",X"A7",X"C8",X"1C",X"E6",X"C8",X"1E",
		X"C1",X"02",X"10",X"24",X"02",X"31",X"BD",X"64",X"39",X"86",X"01",X"BD",X"D6",X"BA",X"6A",X"C8",
		X"1C",X"26",X"EA",X"6A",X"C8",X"1D",X"26",X"DD",X"A6",X"4C",X"26",X"0A",X"86",X"06",X"8D",X"59",
		X"B6",X"99",X"0A",X"A7",X"C8",X"21",X"EC",X"C8",X"11",X"47",X"56",X"ED",X"4D",X"EC",X"C8",X"13",
		X"47",X"56",X"ED",X"4F",X"E6",X"C8",X"1E",X"C1",X"02",X"10",X"24",X"01",X"FA",X"BD",X"64",X"39",
		X"A6",X"4C",X"27",X"29",X"10",X"AE",X"06",X"2A",X"09",X"10",X"AE",X"2A",X"10",X"AC",X"C8",X"17",
		X"6F",X"06",X"10",X"AE",X"C8",X"17",X"EC",X"35",X"A3",X"4A",X"26",X"03",X"BD",X"64",X"25",X"6F",
		X"4C",X"33",X"A4",X"BD",X"6B",X"F3",X"25",X"05",X"86",X"2D",X"BD",X"D6",X"BA",X"AE",X"47",X"6F",
		X"06",X"86",X"03",X"8E",X"61",X"DA",X"7E",X"D6",X"BC",X"A7",X"C8",X"15",X"35",X"06",X"ED",X"C8",
		X"1F",X"AE",X"47",X"6C",X"02",X"E6",X"C8",X"1E",X"C1",X"02",X"10",X"24",X"01",X"A9",X"1A",X"50",
		X"AE",X"47",X"10",X"AE",X"1A",X"10",X"BF",X"CA",X"02",X"EC",X"3E",X"FD",X"CA",X"06",X"A6",X"11",
		X"27",X"2D",X"E6",X"13",X"FD",X"CA",X"04",X"C6",X"0A",X"A6",X"C8",X"15",X"85",X"01",X"26",X"07",
		X"86",X"22",X"B7",X"CA",X"01",X"C6",X"1A",X"A6",X"12",X"2A",X"02",X"CA",X"20",X"F7",X"CA",X"00",
		X"6A",X"C8",X"15",X"27",X"0A",X"1C",X"AF",X"86",X"03",X"8E",X"62",X"F5",X"7E",X"D6",X"BC",X"1C",
		X"AF",X"6F",X"02",X"86",X"03",X"BD",X"D6",X"BA",X"6E",X"D8",X"1F",X"67",X"4D",X"66",X"4E",X"67",
		X"4F",X"66",X"C8",X"10",X"39",X"A6",X"39",X"81",X"0C",X"23",X"79",X"34",X"20",X"10",X"8E",X"99",
		X"0C",X"8C",X"99",X"91",X"27",X"04",X"10",X"8E",X"99",X"15",X"33",X"84",X"BD",X"6B",X"F3",X"DE",
		X"1C",X"24",X"11",X"EC",X"4D",X"ED",X"C8",X"11",X"EC",X"4F",X"ED",X"C8",X"13",X"86",X"01",X"A7",
		X"4C",X"7E",X"62",X"5E",X"A6",X"25",X"2F",X"1E",X"8B",X"99",X"19",X"A7",X"25",X"6C",X"24",X"31",
		X"84",X"BD",X"D6",X"8B",X"8D",X"52",X"33",X"10",X"AF",X"0B",X"4F",X"5F",X"35",X"40",X"A7",X"46",
		X"ED",X"27",X"ED",X"31",X"20",X"02",X"31",X"84",X"C6",X"03",X"BD",X"D6",X"8B",X"5E",X"8B",X"03",
		X"10",X"AF",X"07",X"5A",X"26",X"F4",X"DE",X"1C",X"86",X"0A",X"A7",X"C8",X"1B",X"AE",X"47",X"10",
		X"AE",X"4A",X"BD",X"64",X"70",X"6A",X"C8",X"1B",X"10",X"27",X"FE",X"E8",X"86",X"01",X"8E",X"63",
		X"BD",X"7E",X"D6",X"BC",X"BD",X"64",X"39",X"6A",X"C8",X"1A",X"26",X"41",X"86",X"02",X"A7",X"C8",
		X"1A",X"A6",X"05",X"4C",X"81",X"03",X"25",X"15",X"8E",X"E6",X"6A",X"BD",X"E6",X"AA",X"AE",X"47",
		X"A6",X"C8",X"19",X"27",X"08",X"86",X"02",X"BD",X"62",X"E9",X"AE",X"47",X"4F",X"1A",X"50",X"E6",
		X"11",X"10",X"27",X"00",X"C2",X"A7",X"05",X"10",X"AE",X"08",X"C6",X"05",X"3D",X"31",X"A5",X"EC",
		X"15",X"E3",X"22",X"ED",X"15",X"A6",X"17",X"AB",X"24",X"A7",X"17",X"1C",X"AF",X"86",X"03",X"8E",
		X"61",X"DA",X"7E",X"D6",X"BC",X"34",X"10",X"BE",X"99",X"CE",X"EC",X"4A",X"10",X"B3",X"99",X"86",
		X"27",X"03",X"BE",X"99",X"86",X"AF",X"4A",X"35",X"90",X"A6",X"4F",X"2A",X"01",X"40",X"81",X"0C",
		X"23",X"01",X"3F",X"AE",X"47",X"10",X"AE",X"4A",X"A6",X"31",X"27",X"09",X"EE",X"2A",X"BD",X"6B",
		X"F3",X"DE",X"1C",X"24",X"05",X"8D",X"CE",X"10",X"AE",X"4A",X"A6",X"11",X"27",X"69",X"D6",X"D1",
		X"27",X"0E",X"81",X"49",X"CC",X"FF",X"00",X"25",X"03",X"CC",X"01",X"00",X"E3",X"15",X"20",X"19",
		X"EC",X"15",X"10",X"A3",X"35",X"24",X"04",X"E3",X"4D",X"E3",X"4D",X"A3",X"4D",X"81",X"08",X"24",
		X"02",X"86",X"08",X"81",X"7F",X"25",X"02",X"86",X"7F",X"ED",X"15",X"EC",X"17",X"10",X"A3",X"37",
		X"24",X"04",X"E3",X"4F",X"E3",X"4F",X"A3",X"4F",X"81",X"41",X"24",X"02",X"86",X"41",X"81",X"C9",
		X"25",X"02",X"86",X"C9",X"ED",X"17",X"39",X"10",X"AE",X"47",X"8E",X"8F",X"48",X"86",X"32",X"BD",
		X"D6",X"76",X"A6",X"31",X"E6",X"33",X"C3",X"06",X"0A",X"ED",X"88",X"28",X"86",X"FF",X"A7",X"23",
		X"86",X"03",X"BD",X"D6",X"BA",X"AE",X"47",X"9C",X"77",X"26",X"04",X"0F",X"77",X"20",X"02",X"0F",
		X"79",X"1C",X"AF",X"BD",X"D7",X"84",X"BD",X"DC",X"73",X"0A",X"76",X"7E",X"D6",X"C5",X"00",X"FF",
		X"00",X"FF",X"00",X"80",X"00",X"00",X"86",X"42",X"32",X"23",X"22",X"E0",X"00",X"FF",X"00",X"FF",
		X"00",X"80",X"00",X"00",X"86",X"42",X"33",X"33",X"22",X"E8",X"00",X"C0",X"00",X"80",X"00",X"20",
		X"00",X"00",X"43",X"21",X"32",X"12",X"11",X"E0",X"00",X"40",X"00",X"30",X"00",X"20",X"00",X"10",
		X"86",X"42",X"33",X"33",X"22",X"F8",X"00",X"40",X"00",X"30",X"00",X"20",X"00",X"10",X"86",X"42",
		X"33",X"33",X"22",X"F0",X"00",X"40",X"00",X"30",X"00",X"1E",X"00",X"00",X"64",X"21",X"33",X"22",
		X"22",X"FB",X"00",X"03",X"00",X"02",X"00",X"02",X"00",X"00",X"86",X"42",X"43",X"23",X"21",X"FF",
		X"04",X"80",X"02",X"80",X"02",X"00",X"02",X"00",X"53",X"21",X"32",X"22",X"22",X"B0",X"01",X"40",
		X"01",X"D0",X"01",X"C0",X"02",X"30",X"FA",X"52",X"A5",X"35",X"32",X"15",X"02",X"80",X"03",X"00",
		X"03",X"C0",X"03",X"C0",X"FA",X"52",X"A5",X"35",X"32",X"30",X"00",X"F0",X"00",X"80",X"00",X"30",
		X"00",X"06",X"44",X"32",X"54",X"35",X"32",X"FB",X"01",X"40",X"01",X"80",X"02",X"00",X"03",X"80",
		X"44",X"32",X"54",X"35",X"32",X"40",X"00",X"01",X"00",X"02",X"00",X"02",X"00",X"05",X"75",X"44",
		X"54",X"34",X"53",X"01",X"00",X"90",X"00",X"80",X"00",X"72",X"00",X"45",X"44",X"32",X"43",X"34",
		X"32",X"FD",X"00",X"70",X"00",X"64",X"00",X"50",X"00",X"15",X"44",X"32",X"43",X"34",X"32",X"F6",
		X"00",X"0E",X"00",X"0C",X"00",X"0A",X"00",X"06",X"44",X"32",X"33",X"34",X"32",X"FF",X"00",X"40",
		X"00",X"45",X"00",X"50",X"00",X"70",X"32",X"21",X"21",X"11",X"21",X"05",X"00",X"A0",X"00",X"80",
		X"00",X"70",X"00",X"40",X"44",X"33",X"43",X"32",X"21",X"E0",X"00",X"FF",X"00",X"E0",X"00",X"C0",
		X"00",X"90",X"87",X"66",X"76",X"54",X"42",X"C0",X"96",X"39",X"48",X"2B",X"08",X"81",X"06",X"27",
		X"07",X"D6",X"8D",X"26",X"61",X"6E",X"D8",X"07",X"4F",X"5F",X"FD",X"99",X"82",X"FD",X"99",X"CA",
		X"FD",X"BF",X"2A",X"FD",X"BF",X"2C",X"FD",X"BF",X"2E",X"FD",X"BF",X"30",X"97",X"68",X"10",X"8E",
		X"40",X"A0",X"BD",X"69",X"56",X"8E",X"E6",X"A4",X"BD",X"E6",X"AA",X"BD",X"D6",X"8B",X"79",X"7B",
		X"24",X"86",X"7D",X"BD",X"D6",X"BA",X"8E",X"37",X"E6",X"86",X"51",X"BD",X"D6",X"76",X"86",X"01",
		X"BD",X"D6",X"BA",X"B6",X"BF",X"35",X"26",X"05",X"86",X"FF",X"BD",X"D6",X"BA",X"0F",X"39",X"BD",
		X"D7",X"0D",X"BD",X"7F",X"0B",X"BD",X"D6",X"8B",X"79",X"7B",X"24",X"8E",X"37",X"E6",X"86",X"51",
		X"BD",X"D6",X"76",X"7E",X"D6",X"C5",X"10",X"8E",X"68",X"0F",X"85",X"02",X"26",X"08",X"F6",X"99",
		X"11",X"27",X"03",X"BD",X"67",X"CB",X"31",X"24",X"96",X"39",X"85",X"02",X"26",X"08",X"F6",X"99",
		X"1A",X"27",X"03",X"BD",X"67",X"CB",X"0C",X"87",X"96",X"87",X"81",X"23",X"23",X"04",X"80",X"06",
		X"20",X"F8",X"BD",X"E7",X"FD",X"C6",X"05",X"BD",X"37",X"B9",X"86",X"C3",X"BD",X"D6",X"BA",X"0F",
		X"8D",X"D6",X"D0",X"F7",X"99",X"04",X"8E",X"CC",X"14",X"BD",X"37",X"BF",X"A7",X"E2",X"8E",X"64",
		X"DE",X"10",X"8E",X"98",X"D3",X"E6",X"22",X"27",X"04",X"6A",X"22",X"26",X"2A",X"E6",X"E4",X"CB",
		X"10",X"57",X"E6",X"85",X"25",X"04",X"54",X"54",X"54",X"54",X"C4",X"0F",X"E7",X"22",X"E6",X"0D",
		X"1D",X"2B",X"09",X"E3",X"A4",X"10",X"A3",X"06",X"2D",X"0B",X"20",X"07",X"E3",X"A4",X"10",X"A3",
		X"06",X"2E",X"02",X"EC",X"06",X"ED",X"A4",X"30",X"0E",X"31",X"23",X"8C",X"65",X"E8",X"25",X"C5",
		X"35",X"02",X"B6",X"99",X"04",X"97",X"D0",X"0F",X"7D",X"0F",X"CB",X"0C",X"85",X"0C",X"68",X"96",
		X"87",X"80",X"06",X"24",X"FC",X"8B",X"06",X"8E",X"68",X"17",X"E6",X"86",X"C4",X"0F",X"D7",X"8E",
		X"E6",X"86",X"C4",X"F0",X"D7",X"8F",X"81",X"04",X"26",X"1F",X"86",X"10",X"97",X"8B",X"0F",X"85",
		X"0C",X"75",X"86",X"90",X"B7",X"99",X"04",X"96",X"87",X"81",X"16",X"24",X"06",X"CC",X"68",X"F3",
		X"7E",X"67",X"AD",X"CC",X"68",X"ED",X"7E",X"67",X"AD",X"81",X"02",X"26",X"28",X"86",X"69",X"B7",
		X"99",X"04",X"86",X"01",X"97",X"83",X"0C",X"86",X"C6",X"2C",X"96",X"87",X"81",X"0C",X"25",X"01",
		X"5F",X"D7",X"BA",X"81",X"12",X"25",X"09",X"0F",X"85",X"0F",X"D1",X"CC",X"68",X"DF",X"20",X"5D",
		X"CC",X"68",X"E3",X"20",X"58",X"4D",X"26",X"1C",X"96",X"8C",X"97",X"8B",X"0F",X"83",X"96",X"87",
		X"81",X"0C",X"24",X"07",X"0C",X"86",X"CC",X"68",X"37",X"20",X"42",X"0F",X"85",X"0F",X"D1",X"CC",
		X"68",X"1D",X"20",X"39",X"81",X"01",X"26",X"05",X"CC",X"68",X"42",X"20",X"30",X"81",X"03",X"26",
		X"1A",X"0F",X"D1",X"0F",X"85",X"86",X"C0",X"B7",X"99",X"04",X"86",X"80",X"D6",X"87",X"C1",X"09",
		X"25",X"02",X"86",X"82",X"97",X"83",X"CC",X"68",X"D3",X"20",X"12",X"0F",X"68",X"0F",X"85",X"0C",
		X"86",X"CC",X"69",X"91",X"DD",X"CE",X"86",X"82",X"97",X"83",X"CC",X"69",X"04",X"ED",X"47",X"86",
		X"19",X"A7",X"4D",X"A7",X"4A",X"8B",X"14",X"A7",X"4B",X"8B",X"23",X"A7",X"4C",X"BD",X"D6",X"8B",
		X"DD",X"3F",X"14",X"86",X"03",X"8E",X"65",X"E8",X"7E",X"D6",X"BC",X"BD",X"D6",X"8B",X"E8",X"E6",
		X"27",X"EE",X"A4",X"EF",X"07",X"EE",X"22",X"EF",X"09",X"86",X"3C",X"A7",X"0B",X"BD",X"D6",X"8B",
		X"E8",X"EB",X"19",X"C5",X"F0",X"26",X"02",X"CA",X"F0",X"E7",X"07",X"EC",X"21",X"ED",X"08",X"A6",
		X"23",X"8B",X"0B",X"C6",X"3C",X"ED",X"0A",X"BD",X"D6",X"8B",X"E8",X"E6",X"27",X"EC",X"A4",X"86",
		X"DF",X"ED",X"07",X"EC",X"22",X"C3",X"0A",X"0B",X"ED",X"09",X"C6",X"3C",X"E7",X"0B",X"39",X"5E",
		X"44",X"2A",X"C0",X"5F",X"22",X"56",X"C0",X"44",X"33",X"77",X"55",X"66",X"22",X"C6",X"01",X"E7",
		X"4A",X"BD",X"69",X"36",X"BD",X"69",X"19",X"86",X"03",X"8E",X"65",X"E8",X"7E",X"D6",X"BC",X"6A",
		X"49",X"26",X"07",X"0C",X"85",X"20",X"03",X"BD",X"68",X"B4",X"86",X"03",X"8E",X"65",X"E8",X"7E",
		X"D6",X"BC",X"96",X"87",X"81",X"07",X"96",X"7D",X"C6",X"01",X"25",X"02",X"8B",X"02",X"81",X"05",
		X"25",X"01",X"5C",X"96",X"87",X"81",X"13",X"25",X"02",X"C6",X"02",X"D1",X"7B",X"23",X"0A",X"0C",
		X"7B",X"8E",X"86",X"1C",X"86",X"26",X"BD",X"D6",X"76",X"86",X"03",X"8E",X"65",X"E8",X"7E",X"D6",
		X"BC",X"A6",X"4B",X"26",X"3B",X"96",X"88",X"26",X"35",X"9E",X"7E",X"2A",X"04",X"E6",X"13",X"2A",
		X"2D",X"BD",X"5D",X"BF",X"8A",X"28",X"C6",X"50",X"3D",X"A7",X"4B",X"BD",X"D6",X"8B",X"81",X"E5",
		X"23",X"BD",X"EA",X"FA",X"2A",X"02",X"86",X"04",X"A7",X"08",X"8E",X"98",X"A3",X"6C",X"86",X"D6",
		X"83",X"2A",X"08",X"BD",X"5D",X"BF",X"C6",X"05",X"3D",X"97",X"84",X"C6",X"01",X"39",X"5F",X"39",
		X"6A",X"4B",X"20",X"FA",X"E6",X"4A",X"26",X"17",X"D6",X"74",X"26",X"11",X"86",X"28",X"A7",X"4A",
		X"86",X"25",X"8E",X"82",X"C8",X"BD",X"D6",X"76",X"0C",X"74",X"0C",X"88",X"39",X"5F",X"39",X"6A",
		X"4A",X"20",X"FA",X"BD",X"68",X"71",X"C6",X"01",X"96",X"87",X"81",X"07",X"25",X"58",X"5C",X"C6",
		X"01",X"8D",X"53",X"8D",X"34",X"86",X"03",X"8E",X"65",X"E8",X"7E",X"D6",X"BC",X"8D",X"2A",X"C6",
		X"03",X"20",X"02",X"C6",X"04",X"D1",X"74",X"23",X"EC",X"E6",X"4A",X"26",X"03",X"BD",X"68",X"BC",
		X"6A",X"4A",X"20",X"E1",X"BD",X"68",X"71",X"27",X"06",X"86",X"32",X"A7",X"4B",X"20",X"D6",X"D6",
		X"87",X"C1",X"0B",X"25",X"D0",X"8D",X"02",X"20",X"CC",X"96",X"7B",X"26",X"18",X"6A",X"4C",X"26",
		X"14",X"BD",X"5D",X"BF",X"8A",X"28",X"C6",X"64",X"3D",X"A7",X"4C",X"0C",X"7B",X"8E",X"86",X"1C",
		X"86",X"26",X"BD",X"D6",X"76",X"39",X"D1",X"76",X"23",X"14",X"0C",X"CB",X"6A",X"4D",X"26",X"0E",
		X"86",X"14",X"A7",X"4D",X"8E",X"60",X"CE",X"86",X"29",X"BD",X"D6",X"76",X"0C",X"76",X"86",X"03",
		X"8E",X"65",X"E8",X"7E",X"D6",X"BC",X"34",X"16",X"C6",X"78",X"20",X"15",X"34",X"16",X"BD",X"D6",
		X"8B",X"E8",X"E6",X"27",X"E7",X"07",X"86",X"44",X"A7",X"08",X"10",X"AF",X"09",X"C6",X"3C",X"E7",
		X"0B",X"BD",X"D6",X"8B",X"E8",X"E6",X"27",X"E7",X"0B",X"CC",X"5C",X"44",X"ED",X"07",X"31",X"A9",
		X"FD",X"F1",X"10",X"AF",X"09",X"35",X"96",X"8E",X"E6",X"6D",X"BD",X"E6",X"AA",X"6E",X"9F",X"98",
		X"CE",X"96",X"87",X"81",X"06",X"25",X"05",X"CC",X"09",X"09",X"DD",X"CC",X"BE",X"9A",X"16",X"AF",
		X"47",X"A6",X"15",X"E6",X"17",X"ED",X"4A",X"86",X"08",X"A7",X"49",X"BE",X"9A",X"38",X"A6",X"11",
		X"10",X"27",X"6D",X"11",X"E6",X"13",X"ED",X"4C",X"6F",X"4E",X"AE",X"47",X"A6",X"11",X"10",X"27",
		X"6D",X"03",X"EC",X"4A",X"A0",X"4C",X"2A",X"01",X"40",X"97",X"3E",X"E0",X"4D",X"2A",X"01",X"50",
		X"57",X"D0",X"3E",X"24",X"13",X"6A",X"4E",X"0F",X"3E",X"A6",X"49",X"8E",X"6A",X"78",X"30",X"86",
		X"EC",X"84",X"6D",X"4E",X"2A",X"02",X"1E",X"89",X"47",X"AB",X"4C",X"A0",X"4A",X"97",X"45",X"2A",
		X"01",X"40",X"48",X"24",X"02",X"86",X"FF",X"EB",X"4D",X"E0",X"4B",X"C0",X"08",X"D7",X"46",X"2A",
		X"01",X"50",X"DD",X"3F",X"6D",X"4E",X"2A",X"28",X"96",X"CC",X"D6",X"3F",X"8D",X"74",X"48",X"48",
		X"D6",X"46",X"2A",X"03",X"50",X"0C",X"3E",X"8D",X"69",X"DD",X"41",X"96",X"CC",X"5F",X"47",X"56",
		X"47",X"56",X"47",X"56",X"0D",X"45",X"2A",X"04",X"43",X"50",X"82",X"FF",X"DD",X"3F",X"20",X"23",
		X"96",X"CD",X"D6",X"40",X"8D",X"4C",X"48",X"48",X"D6",X"45",X"2A",X"03",X"50",X"0C",X"3E",X"8D",
		X"41",X"47",X"56",X"DD",X"3F",X"96",X"CD",X"5F",X"47",X"59",X"47",X"59",X"0D",X"46",X"2A",X"01",
		X"40",X"DD",X"41",X"EC",X"4A",X"CB",X"08",X"DD",X"43",X"CC",X"0C",X"08",X"BD",X"88",X"E4",X"6A",
		X"49",X"6A",X"49",X"10",X"2B",X"6C",X"5E",X"BE",X"9A",X"38",X"A6",X"11",X"10",X"27",X"6C",X"55",
		X"86",X"01",X"8E",X"69",X"D7",X"7E",X"D6",X"BC",X"F6",X"00",X"0A",X"00",X"EC",X"00",X"14",X"00",
		X"00",X"00",X"97",X"3C",X"4F",X"8D",X"14",X"97",X"43",X"1F",X"98",X"5F",X"8D",X"0D",X"1F",X"89",
		X"96",X"43",X"0D",X"3E",X"27",X"04",X"43",X"50",X"82",X"FF",X"39",X"97",X"47",X"86",X"08",X"97",
		X"3D",X"96",X"47",X"58",X"49",X"91",X"3C",X"25",X"03",X"90",X"3C",X"5C",X"0A",X"3D",X"26",X"F3",
		X"1E",X"89",X"39",X"BE",X"9A",X"16",X"AF",X"47",X"86",X"04",X"A7",X"49",X"03",X"BC",X"2B",X"01",
		X"4F",X"A7",X"4A",X"AE",X"47",X"A6",X"11",X"10",X"27",X"6B",X"FA",X"E6",X"17",X"C3",X"01",X"07",
		X"DD",X"43",X"8E",X"6A",X"F9",X"A6",X"4A",X"48",X"48",X"30",X"86",X"EC",X"84",X"DD",X"3F",X"EC",
		X"02",X"DD",X"41",X"CC",X"0C",X"08",X"BD",X"88",X"E4",X"6C",X"4A",X"6A",X"49",X"10",X"27",X"6B",
		X"D4",X"86",X"01",X"8E",X"6A",X"C3",X"7E",X"D6",X"BC",X"00",X"00",X"FD",X"00",X"01",X"80",X"00",
		X"00",X"00",X"00",X"03",X"00",X"FE",X"80",X"00",X"00",X"00",X"C0",X"FE",X"80",X"00",X"C0",X"01",
		X"80",X"FF",X"40",X"01",X"80",X"FF",X"40",X"FE",X"80",X"DE",X"1C",X"AE",X"47",X"10",X"AE",X"0A",
		X"86",X"0F",X"A7",X"4D",X"33",X"A4",X"BD",X"6B",X"F3",X"24",X"0A",X"D6",X"F2",X"E7",X"A8",X"26",
		X"CC",X"74",X"82",X"ED",X"2A",X"DE",X"1C",X"CC",X"FB",X"80",X"ED",X"49",X"ED",X"A8",X"29",X"A6",
		X"13",X"8B",X"14",X"A7",X"4E",X"AE",X"47",X"E6",X"4D",X"2B",X"08",X"6A",X"4D",X"26",X"0A",X"C6",
		X"FC",X"E7",X"03",X"A6",X"17",X"A1",X"4E",X"24",X"0A",X"8D",X"35",X"86",X"01",X"8E",X"6B",X"45",
		X"7E",X"D6",X"BC",X"8D",X"2B",X"8E",X"E6",X"89",X"BD",X"E6",X"AA",X"86",X"07",X"BD",X"D6",X"BA",
		X"AE",X"47",X"10",X"AE",X"0A",X"EC",X"A8",X"29",X"10",X"83",X"02",X"00",X"23",X"0E",X"47",X"56",
		X"47",X"56",X"43",X"50",X"82",X"FF",X"E3",X"A8",X"29",X"ED",X"A8",X"29",X"ED",X"49",X"20",X"C9",
		X"10",X"AE",X"1A",X"EC",X"15",X"E3",X"4B",X"10",X"83",X"06",X"80",X"25",X"15",X"AB",X"3E",X"10",
		X"83",X"8F",X"00",X"22",X"06",X"A0",X"3E",X"ED",X"15",X"20",X"14",X"CC",X"8F",X"00",X"A0",X"3E",
		X"20",X"03",X"CC",X"06",X"80",X"ED",X"15",X"EC",X"4B",X"43",X"50",X"82",X"FF",X"ED",X"4B",X"EC",
		X"49",X"C3",X"00",X"20",X"ED",X"49",X"E3",X"17",X"81",X"3A",X"23",X"13",X"AB",X"3F",X"81",X"D6",
		X"24",X"06",X"A0",X"3F",X"ED",X"17",X"20",X"1A",X"CC",X"D5",X"00",X"A0",X"3F",X"20",X"09",X"A6",
		X"4E",X"80",X"19",X"A7",X"4E",X"CC",X"3B",X"00",X"ED",X"17",X"EC",X"49",X"43",X"50",X"82",X"FF",
		X"ED",X"49",X"39",X"34",X"02",X"96",X"39",X"11",X"83",X"99",X"91",X"27",X"01",X"46",X"46",X"35",
		X"82",X"AE",X"47",X"A6",X"06",X"26",X"36",X"A6",X"11",X"10",X"26",X"02",X"69",X"A6",X"03",X"81",
		X"04",X"26",X"24",X"A6",X"19",X"81",X"08",X"26",X"1E",X"96",X"D1",X"27",X"1A",X"96",X"81",X"81",
		X"02",X"24",X"14",X"0C",X"81",X"31",X"84",X"86",X"30",X"8E",X"89",X"CF",X"BD",X"D6",X"76",X"A6",
		X"35",X"E6",X"37",X"ED",X"07",X"30",X"A4",X"BD",X"D7",X"84",X"7E",X"D6",X"C5",X"10",X"AE",X"06",
		X"A6",X"39",X"85",X"F0",X"26",X"5D",X"EE",X"2A",X"11",X"83",X"9A",X"21",X"23",X"06",X"E6",X"45",
		X"C1",X"22",X"26",X"0A",X"6F",X"06",X"86",X"01",X"8E",X"6C",X"01",X"7E",X"D6",X"BC",X"81",X"0E",
		X"26",X"38",X"A6",X"23",X"81",X"10",X"27",X"32",X"EE",X"2A",X"E6",X"03",X"E7",X"49",X"10",X"8E",
		X"99",X"0C",X"57",X"25",X"07",X"57",X"24",X"22",X"10",X"8E",X"99",X"15",X"A6",X"19",X"44",X"34",
		X"10",X"8E",X"6E",X"AE",X"A6",X"86",X"BD",X"E1",X"2C",X"35",X"10",X"6C",X"C8",X"1E",X"E6",X"C8",
		X"1E",X"C1",X"02",X"25",X"05",X"86",X"20",X"BD",X"E1",X"20",X"BD",X"D7",X"84",X"BD",X"DC",X"73",
		X"7E",X"D6",X"C5",X"85",X"30",X"27",X"37",X"E6",X"45",X"2B",X"A9",X"C6",X"05",X"8E",X"5E",X"96",
		X"85",X"10",X"26",X"05",X"C6",X"10",X"8E",X"5E",X"A0",X"86",X"41",X"BD",X"D6",X"95",X"10",X"AF",
		X"07",X"10",X"AE",X"47",X"10",X"AF",X"09",X"A6",X"23",X"10",X"8E",X"99",X"0C",X"47",X"25",X"07",
		X"47",X"24",X"CD",X"10",X"8E",X"99",X"15",X"1F",X"98",X"BD",X"E1",X"20",X"20",X"C2",X"EE",X"2A",
		X"85",X"80",X"27",X"1E",X"85",X"40",X"26",X"14",X"85",X"01",X"26",X"04",X"E6",X"5B",X"20",X"02",
		X"E6",X"5D",X"26",X"39",X"E6",X"53",X"2A",X"35",X"33",X"A4",X"20",X"19",X"A6",X"53",X"10",X"2A",
		X"FF",X"52",X"E6",X"03",X"C1",X"04",X"26",X"35",X"E6",X"53",X"10",X"2A",X"FF",X"46",X"4F",X"E6",
		X"5B",X"26",X"08",X"EE",X"57",X"BD",X"D5",X"5A",X"7E",X"D6",X"C5",X"E6",X"5D",X"10",X"26",X"FF",
		X"79",X"EE",X"59",X"4C",X"20",X"EF",X"10",X"AE",X"47",X"EE",X"49",X"20",X"17",X"A6",X"03",X"81",
		X"04",X"26",X"0A",X"86",X"02",X"BD",X"D6",X"BA",X"AE",X"47",X"7E",X"6C",X"9A",X"6C",X"02",X"31",
		X"84",X"BD",X"6E",X"0D",X"BD",X"D6",X"8B",X"5E",X"83",X"03",X"10",X"AF",X"09",X"EF",X"07",X"11",
		X"83",X"9A",X"21",X"27",X"5A",X"EC",X"53",X"2A",X"4B",X"1A",X"50",X"AE",X"53",X"6D",X"11",X"10",
		X"27",X"00",X"A5",X"AE",X"5B",X"2A",X"08",X"6F",X"5B",X"BD",X"D7",X"84",X"BD",X"DC",X"73",X"AE",
		X"5D",X"2A",X"08",X"6F",X"5D",X"BD",X"D7",X"84",X"BD",X"DC",X"73",X"9E",X"1C",X"ED",X"07",X"ED",
		X"C8",X"27",X"6F",X"53",X"1C",X"AF",X"CC",X"02",X"80",X"6D",X"3C",X"2B",X"04",X"43",X"50",X"82",
		X"FF",X"ED",X"0B",X"EC",X"51",X"84",X"3F",X"C4",X"FC",X"ED",X"51",X"BD",X"DF",X"C1",X"AF",X"C8",
		X"37",X"7E",X"6B",X"19",X"4F",X"5F",X"ED",X"51",X"9E",X"1C",X"EF",X"0B",X"7E",X"8D",X"52",X"AE",
		X"55",X"E6",X"03",X"2B",X"53",X"1A",X"50",X"E6",X"11",X"27",X"4D",X"31",X"84",X"8E",X"8F",X"48",
		X"86",X"34",X"BD",X"D6",X"76",X"A6",X"31",X"E6",X"33",X"ED",X"88",X"28",X"30",X"A4",X"4F",X"5F",
		X"ED",X"51",X"4A",X"10",X"8E",X"8D",X"37",X"BD",X"8D",X"DD",X"1C",X"AF",X"86",X"02",X"BD",X"D6",
		X"BA",X"CE",X"9A",X"21",X"1A",X"50",X"10",X"8E",X"8D",X"3C",X"BD",X"8D",X"DD",X"86",X"08",X"10",
		X"8E",X"8D",X"37",X"BD",X"8D",X"DD",X"1C",X"AF",X"86",X"5A",X"BD",X"D6",X"BA",X"CE",X"9A",X"21",
		X"86",X"FF",X"A7",X"C8",X"24",X"6F",X"C8",X"23",X"1C",X"AF",X"7E",X"D6",X"C5",X"34",X"36",X"E6",
		X"39",X"54",X"8E",X"E6",X"96",X"BD",X"E6",X"AA",X"8E",X"6E",X"AE",X"A6",X"85",X"E6",X"23",X"11",
		X"83",X"9A",X"21",X"26",X"18",X"10",X"8E",X"99",X"0C",X"54",X"25",X"07",X"54",X"24",X"45",X"10",
		X"8E",X"99",X"15",X"BD",X"E1",X"2C",X"86",X"15",X"BD",X"E1",X"20",X"20",X"37",X"10",X"8E",X"99",
		X"15",X"8E",X"99",X"0C",X"11",X"83",X"99",X"91",X"27",X"07",X"10",X"8E",X"99",X"0C",X"8E",X"99",
		X"15",X"C5",X"03",X"27",X"0C",X"BD",X"E1",X"2C",X"A6",X"53",X"2B",X"18",X"86",X"20",X"BD",X"E1",
		X"20",X"A6",X"53",X"2B",X"0F",X"A6",X"05",X"2F",X"0B",X"8B",X"99",X"19",X"A7",X"05",X"6C",X"04",
		X"9E",X"1C",X"A7",X"0E",X"35",X"B6",X"A6",X"19",X"84",X"0E",X"10",X"8E",X"6E",X"B5",X"31",X"A6",
		X"E6",X"21",X"27",X"22",X"A6",X"49",X"4C",X"A1",X"A4",X"25",X"19",X"A6",X"04",X"5A",X"27",X"0C",
		X"E6",X"4A",X"C4",X"03",X"27",X"06",X"C1",X"03",X"27",X"02",X"4A",X"4A",X"4C",X"84",X"07",X"6C",
		X"4A",X"A7",X"05",X"4F",X"A7",X"49",X"86",X"01",X"8E",X"6C",X"01",X"7E",X"D6",X"BC",X"52",X"52",
		X"04",X"57",X"05",X"52",X"09",X"03",X"01",X"00",X"00",X"06",X"02",X"0C",X"02",X"04",X"01",X"00",
		X"00",X"00",X"00",X"96",X"39",X"2B",X"01",X"39",X"43",X"85",X"03",X"27",X"FA",X"CE",X"99",X"91",
		X"AE",X"55",X"BD",X"6F",X"67",X"A6",X"03",X"81",X"FF",X"27",X"40",X"A6",X"C8",X"23",X"2B",X"05",
		X"BD",X"71",X"A3",X"20",X"36",X"96",X"39",X"85",X"01",X"27",X"0B",X"FC",X"99",X"CE",X"ED",X"C8",
		X"17",X"BD",X"74",X"6E",X"20",X"02",X"DC",X"58",X"6D",X"11",X"27",X"0C",X"AE",X"47",X"27",X"0D",
		X"84",X"F0",X"AA",X"80",X"6D",X"84",X"26",X"03",X"8E",X"00",X"00",X"AF",X"47",X"AE",X"55",X"B4",
		X"99",X"82",X"F4",X"99",X"83",X"BD",X"70",X"22",X"BD",X"E3",X"8D",X"CE",X"99",X"D9",X"AE",X"55",
		X"8D",X"45",X"A6",X"03",X"81",X"FF",X"27",X"3E",X"A6",X"C8",X"23",X"2B",X"03",X"7E",X"71",X"A3",
		X"96",X"39",X"85",X"02",X"27",X"0B",X"FC",X"99",X"86",X"ED",X"C8",X"17",X"BD",X"74",X"6E",X"20",
		X"02",X"DC",X"5C",X"6D",X"11",X"27",X"0C",X"AE",X"47",X"27",X"0D",X"84",X"F0",X"AA",X"80",X"6D",
		X"84",X"26",X"03",X"8E",X"00",X"00",X"AF",X"47",X"AE",X"55",X"B4",X"99",X"CA",X"F4",X"99",X"CB",
		X"BD",X"70",X"22",X"7E",X"E3",X"8D",X"39",X"34",X"76",X"AE",X"5B",X"2A",X"40",X"10",X"AE",X"06",
		X"2A",X"3B",X"EE",X"2A",X"11",X"83",X"D4",X"38",X"27",X"06",X"A6",X"45",X"81",X"22",X"26",X"04",
		X"6F",X"06",X"20",X"29",X"EE",X"66",X"A6",X"39",X"81",X"C0",X"27",X"F4",X"6F",X"5B",X"A6",X"39",
		X"2A",X"19",X"EE",X"2A",X"E6",X"53",X"2A",X"13",X"85",X"01",X"26",X"04",X"EE",X"5B",X"20",X"02",
		X"EE",X"5D",X"2B",X"07",X"33",X"A4",X"BD",X"D5",X"5A",X"20",X"02",X"8D",X"48",X"EE",X"66",X"AE",
		X"5D",X"2A",X"40",X"10",X"AE",X"06",X"2A",X"3B",X"EE",X"2A",X"11",X"83",X"D4",X"38",X"27",X"06",
		X"A6",X"45",X"81",X"22",X"26",X"04",X"6F",X"06",X"20",X"29",X"EE",X"66",X"A6",X"39",X"81",X"C0",
		X"27",X"F4",X"6F",X"5D",X"A6",X"39",X"2A",X"19",X"EE",X"2A",X"E6",X"53",X"2A",X"13",X"85",X"01",
		X"26",X"04",X"EE",X"5B",X"20",X"02",X"EE",X"5D",X"2B",X"07",X"33",X"A4",X"BD",X"D5",X"5A",X"20",
		X"02",X"8D",X"02",X"35",X"F6",X"6C",X"02",X"BD",X"DC",X"73",X"85",X"C0",X"26",X"10",X"EE",X"68",
		X"E6",X"C8",X"2B",X"26",X"05",X"AF",X"C8",X"2B",X"20",X"03",X"AF",X"C8",X"2D",X"39",X"EE",X"2A",
		X"E6",X"C8",X"33",X"26",X"05",X"AF",X"C8",X"33",X"20",X"03",X"AF",X"C8",X"35",X"31",X"84",X"7E",
		X"6E",X"0D",X"34",X"06",X"85",X"01",X"27",X"41",X"EC",X"17",X"A3",X"45",X"81",X"41",X"10",X"25",
		X"00",X"82",X"ED",X"17",X"10",X"AE",X"57",X"EC",X"37",X"A3",X"45",X"ED",X"37",X"10",X"AE",X"59",
		X"EC",X"37",X"A3",X"45",X"ED",X"37",X"10",X"AE",X"53",X"2A",X"06",X"EC",X"37",X"A3",X"45",X"ED",
		X"37",X"10",X"AE",X"5B",X"2A",X"06",X"EC",X"37",X"A3",X"45",X"ED",X"37",X"10",X"AE",X"5D",X"2A",
		X"53",X"EC",X"37",X"A3",X"45",X"ED",X"37",X"20",X"4B",X"85",X"02",X"27",X"47",X"EC",X"17",X"E3",
		X"45",X"11",X"83",X"99",X"D9",X"23",X"04",X"81",X"CC",X"22",X"39",X"81",X"D6",X"22",X"35",X"ED",
		X"17",X"10",X"AE",X"57",X"EC",X"37",X"E3",X"45",X"ED",X"37",X"10",X"AE",X"59",X"EC",X"37",X"E3",
		X"45",X"ED",X"37",X"10",X"AE",X"53",X"2A",X"06",X"EC",X"37",X"E3",X"45",X"ED",X"37",X"10",X"AE",
		X"5B",X"2A",X"06",X"EC",X"37",X"E3",X"45",X"ED",X"37",X"10",X"AE",X"5D",X"2A",X"06",X"EC",X"37",
		X"E3",X"45",X"ED",X"37",X"A6",X"E4",X"85",X"04",X"27",X"43",X"EC",X"15",X"A3",X"43",X"81",X"0F",
		X"10",X"25",X"00",X"91",X"6F",X"C4",X"ED",X"15",X"10",X"AE",X"57",X"EC",X"35",X"A3",X"43",X"ED",
		X"35",X"10",X"AE",X"59",X"EC",X"35",X"A3",X"43",X"ED",X"35",X"10",X"AE",X"53",X"2A",X"06",X"EC",
		X"35",X"A3",X"43",X"ED",X"35",X"10",X"AE",X"5B",X"2A",X"06",X"EC",X"35",X"A3",X"43",X"ED",X"35",
		X"10",X"AE",X"5D",X"2A",X"4D",X"EC",X"35",X"A3",X"43",X"ED",X"35",X"20",X"45",X"85",X"08",X"27",
		X"41",X"EC",X"15",X"E3",X"43",X"81",X"80",X"22",X"4F",X"ED",X"15",X"86",X"01",X"A7",X"C4",X"10",
		X"AE",X"57",X"EC",X"35",X"E3",X"43",X"ED",X"35",X"10",X"AE",X"59",X"EC",X"35",X"E3",X"43",X"ED",
		X"35",X"10",X"AE",X"53",X"2A",X"06",X"EC",X"35",X"E3",X"43",X"ED",X"35",X"10",X"AE",X"5B",X"2A",
		X"06",X"EC",X"35",X"E3",X"43",X"ED",X"35",X"10",X"AE",X"5D",X"2A",X"06",X"EC",X"35",X"E3",X"43",
		X"ED",X"35",X"E6",X"17",X"57",X"E8",X"15",X"C5",X"04",X"26",X"04",X"6F",X"05",X"20",X"04",X"86",
		X"01",X"A7",X"05",X"35",X"86",X"5F",X"20",X"02",X"C6",X"03",X"A6",X"17",X"81",X"8B",X"25",X"05",
		X"B0",X"EA",X"E8",X"20",X"05",X"C8",X"01",X"B0",X"EA",X"EB",X"22",X"01",X"40",X"81",X"0B",X"22",
		X"D1",X"96",X"39",X"11",X"83",X"99",X"D9",X"22",X"C9",X"26",X"06",X"85",X"02",X"27",X"05",X"20",
		X"C1",X"44",X"25",X"BE",X"10",X"AE",X"5D",X"2A",X"08",X"A6",X"39",X"84",X"0E",X"81",X"0A",X"27",
		X"0D",X"10",X"AE",X"5B",X"2A",X"AC",X"A6",X"39",X"84",X"0E",X"81",X"0A",X"26",X"A4",X"E7",X"C8",
		X"23",X"20",X"9F",X"34",X"01",X"1A",X"F0",X"E6",X"C8",X"24",X"C1",X"01",X"10",X"27",X"00",X"58",
		X"10",X"22",X"00",X"94",X"E6",X"47",X"26",X"39",X"10",X"8E",X"71",X"DB",X"BD",X"8D",X"DD",X"AE",
		X"5D",X"AF",X"C8",X"1E",X"AE",X"5B",X"AF",X"C8",X"1C",X"6C",X"C8",X"24",X"10",X"8E",X"71",X"FB",
		X"BD",X"8D",X"DD",X"96",X"8A",X"4C",X"A7",X"C8",X"20",X"35",X"81",X"2A",X"2A",X"E6",X"11",X"27",
		X"0E",X"E6",X"03",X"C1",X"FF",X"27",X"08",X"E6",X"02",X"26",X"04",X"E6",X"06",X"27",X"18",X"32",
		X"64",X"6F",X"C8",X"24",X"C6",X"FF",X"E7",X"C8",X"23",X"35",X"81",X"2A",X"0A",X"EC",X"11",X"ED",
		X"15",X"E6",X"13",X"E7",X"17",X"6F",X"11",X"39",X"E6",X"03",X"C1",X"FF",X"27",X"E3",X"8D",X"12",
		X"A6",X"C8",X"20",X"90",X"8A",X"2A",X"77",X"6C",X"C8",X"24",X"A6",X"C8",X"23",X"BD",X"E9",X"72",
		X"35",X"81",X"AE",X"5D",X"8D",X"1B",X"AC",X"C8",X"1E",X"27",X"05",X"AF",X"C8",X"1E",X"8D",X"0C",
		X"AE",X"5B",X"8D",X"0D",X"AC",X"C8",X"1C",X"27",X"0E",X"AF",X"C8",X"1C",X"30",X"84",X"7E",X"71",
		X"FB",X"2A",X"04",X"A6",X"06",X"26",X"F5",X"39",X"C1",X"20",X"27",X"44",X"24",X"47",X"86",X"FF",
		X"E6",X"C8",X"23",X"C5",X"02",X"27",X"1C",X"40",X"AE",X"5D",X"8D",X"14",X"AE",X"59",X"8D",X"10",
		X"AE",X"55",X"8D",X"0C",X"AE",X"53",X"8D",X"08",X"AE",X"57",X"8D",X"04",X"AE",X"5B",X"20",X"19",
		X"7E",X"5D",X"DB",X"AE",X"57",X"8D",X"F9",X"AE",X"5B",X"8D",X"F5",X"AE",X"55",X"8D",X"F1",X"AE",
		X"53",X"8D",X"ED",X"AE",X"5D",X"8D",X"E9",X"AE",X"59",X"8D",X"E5",X"6C",X"C8",X"24",X"35",X"81",
		X"C6",X"3E",X"E7",X"C8",X"24",X"C1",X"3E",X"25",X"F2",X"C1",X"3F",X"10",X"24",X"00",X"9F",X"6C",
		X"C8",X"24",X"6F",X"5F",X"96",X"39",X"11",X"83",X"99",X"D9",X"22",X"62",X"26",X"3C",X"85",X"02",
		X"27",X"3F",X"96",X"85",X"26",X"05",X"6A",X"C8",X"24",X"35",X"81",X"10",X"BE",X"99",X"86",X"11",
		X"83",X"99",X"D9",X"27",X"04",X"10",X"BE",X"99",X"CE",X"BD",X"5D",X"BF",X"84",X"01",X"E6",X"35",
		X"C1",X"38",X"22",X"02",X"8B",X"02",X"A7",X"C8",X"23",X"BD",X"E9",X"72",X"10",X"AE",X"5D",X"8D",
		X"32",X"25",X"05",X"10",X"AE",X"5B",X"8D",X"2B",X"35",X"81",X"44",X"25",X"C5",X"D6",X"58",X"20",
		X"02",X"D6",X"5C",X"A6",X"C8",X"23",X"88",X"03",X"C5",X"04",X"27",X"06",X"85",X"02",X"26",X"02",
		X"88",X"03",X"C5",X"08",X"27",X"D0",X"85",X"02",X"27",X"CC",X"88",X"03",X"20",X"C8",X"63",X"C8",
		X"24",X"35",X"81",X"34",X"10",X"2A",X"23",X"A6",X"39",X"84",X"0E",X"81",X"0A",X"26",X"1B",X"A6",
		X"39",X"84",X"F1",X"8A",X"06",X"A7",X"39",X"8E",X"00",X"00",X"48",X"AE",X"86",X"AF",X"28",X"EC",
		X"84",X"C3",X"00",X"02",X"ED",X"3A",X"1A",X"01",X"35",X"90",X"1C",X"FE",X"35",X"90",X"6C",X"C8",
		X"24",X"C1",X"5D",X"25",X"2E",X"A6",X"C8",X"23",X"C6",X"03",X"3D",X"10",X"8E",X"EA",X"F1",X"31",
		X"A5",X"A6",X"35",X"E6",X"37",X"8D",X"1E",X"CC",X"FF",X"FF",X"6D",X"53",X"2A",X"02",X"ED",X"51",
		X"A7",X"C8",X"22",X"A7",X"C8",X"23",X"6F",X"C8",X"24",X"BD",X"6B",X"F3",X"24",X"05",X"CC",X"74",
		X"AF",X"ED",X"4A",X"35",X"81",X"34",X"07",X"1A",X"50",X"E6",X"C8",X"25",X"10",X"8E",X"7A",X"9F",
		X"86",X"10",X"3D",X"31",X"A5",X"AE",X"55",X"EC",X"22",X"ED",X"08",X"EC",X"61",X"E7",X"13",X"E7",
		X"17",X"5F",X"E7",X"18",X"E7",X"04",X"E7",X"05",X"E7",X"02",X"ED",X"11",X"ED",X"15",X"BD",X"D8",
		X"C6",X"AE",X"53",X"2A",X"17",X"34",X"40",X"EE",X"55",X"EE",X"48",X"EC",X"47",X"AB",X"63",X"ED",
		X"15",X"ED",X"11",X"A6",X"49",X"AB",X"64",X"BD",X"7C",X"BC",X"35",X"40",X"AE",X"57",X"EC",X"2A",
		X"ED",X"08",X"EC",X"61",X"BD",X"7C",X"C0",X"AE",X"59",X"EC",X"2E",X"ED",X"08",X"EC",X"61",X"BD",
		X"7C",X"C0",X"AE",X"59",X"10",X"AE",X"5D",X"8D",X"24",X"AE",X"57",X"10",X"AE",X"5B",X"8D",X"1D",
		X"6F",X"5F",X"96",X"39",X"85",X"40",X"26",X"09",X"A6",X"53",X"2A",X"05",X"CC",X"FF",X"FF",X"ED",
		X"51",X"CC",X"02",X"00",X"ED",X"45",X"CC",X"01",X"00",X"ED",X"43",X"35",X"87",X"34",X"50",X"2A",
		X"12",X"BD",X"D8",X"D8",X"A6",X"37",X"A7",X"33",X"EC",X"35",X"ED",X"31",X"1F",X"21",X"BD",X"D8",
		X"C6",X"6F",X"02",X"35",X"D0",X"6F",X"C8",X"1A",X"6F",X"C8",X"1B",X"C6",X"FF",X"96",X"39",X"85",
		X"40",X"26",X"04",X"86",X"FF",X"ED",X"51",X"E7",X"C8",X"23",X"CC",X"74",X"47",X"0D",X"23",X"26",
		X"13",X"CC",X"74",X"AF",X"11",X"83",X"99",X"D9",X"26",X"0A",X"86",X"20",X"A7",X"C8",X"24",X"6F",
		X"C8",X"23",X"86",X"74",X"ED",X"4A",X"39",X"C6",X"03",X"E7",X"C8",X"25",X"10",X"8E",X"7A",X"9F",
		X"86",X"10",X"3D",X"31",X"A5",X"AE",X"53",X"EC",X"26",X"ED",X"08",X"4F",X"5F",X"BD",X"7C",X"C0",
		X"6C",X"02",X"AE",X"E4",X"CC",X"74",X"AF",X"ED",X"4A",X"4F",X"5F",X"7E",X"79",X"70",X"EC",X"C8",
		X"1A",X"C1",X"10",X"24",X"08",X"CB",X"10",X"E7",X"C8",X"1B",X"C4",X"03",X"39",X"34",X"50",X"6E",
		X"D8",X"0A",X"6A",X"C8",X"26",X"26",X"E2",X"CC",X"74",X"8C",X"ED",X"4A",X"10",X"AE",X"C8",X"27",
		X"C6",X"03",X"BD",X"ED",X"78",X"7E",X"79",X"70",X"6D",X"5B",X"2A",X"07",X"6D",X"5D",X"2A",X"07",
		X"1A",X"01",X"39",X"6D",X"5D",X"2A",X"05",X"6D",X"C8",X"15",X"26",X"F4",X"1C",X"FE",X"39",X"BD",
		X"5D",X"BF",X"A7",X"C8",X"13",X"BD",X"5D",X"BF",X"A7",X"C8",X"14",X"6F",X"C8",X"15",X"BD",X"5D",
		X"BF",X"91",X"DA",X"22",X"03",X"63",X"C8",X"15",X"6F",X"C8",X"12",X"8D",X"CB",X"24",X"0A",X"CC",
		X"77",X"AD",X"ED",X"4A",X"4F",X"5F",X"7E",X"79",X"70",X"10",X"AE",X"C8",X"17",X"A6",X"35",X"E6",
		X"4E",X"27",X"06",X"81",X"3E",X"22",X"06",X"20",X"10",X"81",X"56",X"22",X"04",X"E6",X"4E",X"27",
		X"0A",X"A7",X"4E",X"10",X"8E",X"76",X"14",X"20",X"06",X"6F",X"4E",X"10",X"8E",X"75",X"08",X"10",
		X"AF",X"4A",X"86",X"3C",X"A7",X"4F",X"6E",X"A4",X"A6",X"53",X"2A",X"06",X"96",X"85",X"10",X"27",
		X"77",X"AD",X"6A",X"4F",X"10",X"27",X"FF",X"97",X"A6",X"4F",X"84",X"01",X"27",X"09",X"7E",X"75",
		X"F0",X"6A",X"4F",X"10",X"27",X"FF",X"88",X"10",X"9E",X"7E",X"10",X"27",X"00",X"BD",X"A6",X"35",
		X"81",X"6F",X"27",X"12",X"81",X"1D",X"10",X"27",X"00",X"B1",X"34",X"10",X"AE",X"2A",X"A6",X"0D",
		X"35",X"10",X"10",X"2F",X"00",X"A5",X"CC",X"75",X"21",X"ED",X"4A",X"4F",X"E6",X"14",X"CB",X"02",
		X"E0",X"37",X"27",X"10",X"22",X"53",X"5C",X"27",X"0B",X"5C",X"27",X"08",X"5C",X"27",X"05",X"5C",
		X"27",X"02",X"86",X"02",X"E6",X"15",X"C4",X"FE",X"C1",X"70",X"25",X"0E",X"C1",X"76",X"27",X"16",
		X"22",X"04",X"8A",X"08",X"20",X"10",X"8A",X"04",X"20",X"0C",X"C1",X"68",X"27",X"08",X"22",X"04",
		X"8A",X"08",X"20",X"02",X"8A",X"04",X"4D",X"26",X"10",X"E6",X"35",X"C1",X"6F",X"26",X"0A",X"E6",
		X"5B",X"26",X"3E",X"E6",X"5D",X"26",X"3A",X"20",X"0C",X"E6",X"5B",X"10",X"26",X"03",X"15",X"E6",
		X"5D",X"10",X"26",X"03",X"0F",X"5F",X"7E",X"79",X"70",X"A6",X"5B",X"10",X"26",X"03",X"05",X"A6",
		X"5D",X"10",X"26",X"02",X"FF",X"E6",X"35",X"CB",X"01",X"86",X"09",X"E1",X"15",X"25",X"E6",X"86",
		X"05",X"C0",X"11",X"E1",X"15",X"25",X"DE",X"26",X"04",X"86",X"01",X"20",X"D8",X"86",X"09",X"20",
		X"D4",X"CC",X"79",X"49",X"ED",X"4A",X"E6",X"35",X"CB",X"01",X"E1",X"15",X"24",X"05",X"CC",X"80",
		X"01",X"20",X"03",X"CC",X"80",X"02",X"ED",X"4C",X"7E",X"79",X"70",X"CC",X"75",X"08",X"ED",X"4A",
		X"A6",X"15",X"84",X"FE",X"6D",X"5D",X"2A",X"0A",X"81",X"76",X"10",X"27",X"01",X"1C",X"25",X"0A",
		X"20",X"0D",X"81",X"68",X"10",X"27",X"01",X"12",X"22",X"05",X"86",X"08",X"7E",X"77",X"1B",X"86",
		X"04",X"7E",X"77",X"1B",X"A6",X"53",X"2A",X"06",X"96",X"85",X"10",X"27",X"76",X"A1",X"6A",X"4F",
		X"10",X"27",X"FE",X"8B",X"A6",X"4F",X"84",X"01",X"27",X"09",X"7E",X"76",X"FC",X"6A",X"4F",X"10",
		X"27",X"FE",X"7C",X"10",X"9E",X"7E",X"10",X"27",X"00",X"BD",X"A6",X"35",X"81",X"1D",X"27",X"12",
		X"81",X"6F",X"10",X"27",X"00",X"B1",X"34",X"10",X"AE",X"2A",X"A6",X"0D",X"35",X"10",X"10",X"2C",
		X"00",X"A5",X"CC",X"76",X"2D",X"ED",X"4A",X"4F",X"E6",X"14",X"CB",X"02",X"E0",X"37",X"27",X"10",
		X"22",X"53",X"5C",X"27",X"0B",X"5C",X"27",X"08",X"5C",X"27",X"05",X"5C",X"27",X"02",X"86",X"02",
		X"E6",X"15",X"C4",X"FE",X"C1",X"1E",X"22",X"0E",X"C1",X"16",X"27",X"16",X"22",X"04",X"8A",X"08",
		X"20",X"10",X"8A",X"04",X"20",X"0C",X"C1",X"24",X"27",X"08",X"22",X"04",X"8A",X"08",X"20",X"02",
		X"8A",X"04",X"4D",X"26",X"10",X"E6",X"35",X"C1",X"1D",X"26",X"0A",X"E6",X"5B",X"26",X"3E",X"E6",
		X"5D",X"26",X"3A",X"20",X"0C",X"E6",X"5B",X"10",X"26",X"02",X"09",X"E6",X"5D",X"10",X"26",X"02",
		X"03",X"5F",X"7E",X"79",X"70",X"A6",X"5B",X"10",X"26",X"01",X"F9",X"A6",X"5D",X"10",X"26",X"01",
		X"F3",X"E6",X"35",X"CB",X"01",X"86",X"05",X"E1",X"15",X"22",X"E6",X"86",X"09",X"C0",X"EE",X"E1",
		X"15",X"22",X"DE",X"26",X"04",X"86",X"01",X"20",X"D8",X"86",X"05",X"20",X"D4",X"CC",X"79",X"49",
		X"ED",X"4A",X"E6",X"35",X"CB",X"01",X"E1",X"15",X"24",X"05",X"CC",X"80",X"01",X"20",X"03",X"CC",
		X"80",X"02",X"ED",X"4C",X"7E",X"79",X"70",X"CC",X"76",X"14",X"ED",X"4A",X"A6",X"15",X"84",X"FE",
		X"6D",X"5B",X"2A",X"08",X"81",X"16",X"27",X"12",X"22",X"08",X"20",X"0A",X"81",X"24",X"27",X"0A",
		X"25",X"04",X"86",X"04",X"20",X"05",X"86",X"08",X"20",X"01",X"4F",X"5F",X"BD",X"74",X"98",X"10",
		X"25",X"00",X"8A",X"34",X"06",X"A6",X"C8",X"13",X"91",X"D4",X"25",X"34",X"10",X"AE",X"C8",X"17",
		X"E6",X"37",X"CB",X"05",X"E0",X"17",X"24",X"09",X"50",X"C1",X"63",X"25",X"0C",X"86",X"01",X"20",
		X"3F",X"C1",X"63",X"25",X"04",X"86",X"02",X"20",X"37",X"54",X"C1",X"0A",X"23",X"17",X"A6",X"35",
		X"A0",X"15",X"24",X"01",X"40",X"34",X"04",X"A0",X"E0",X"24",X"01",X"40",X"81",X"0F",X"23",X"29",
		X"35",X"06",X"7E",X"79",X"70",X"E6",X"17",X"C1",X"D4",X"22",X"13",X"C1",X"43",X"22",X"04",X"86",
		X"02",X"20",X"0D",X"A6",X"C8",X"12",X"26",X"08",X"86",X"02",X"E0",X"37",X"22",X"02",X"86",X"01",
		X"A7",X"C8",X"12",X"AA",X"E4",X"A7",X"E4",X"20",X"D7",X"E6",X"17",X"C1",X"D4",X"22",X"13",X"C1",
		X"43",X"22",X"04",X"86",X"02",X"20",X"0D",X"A6",X"C8",X"12",X"26",X"08",X"86",X"02",X"E0",X"37",
		X"25",X"02",X"86",X"01",X"A7",X"C8",X"12",X"AA",X"E4",X"A7",X"E4",X"20",X"B3",X"10",X"AE",X"C8",
		X"17",X"BD",X"5D",X"BF",X"D6",X"E0",X"58",X"3D",X"1F",X"89",X"4F",X"D0",X"E0",X"82",X"00",X"EB",
		X"37",X"89",X"00",X"2B",X"06",X"10",X"83",X"00",X"43",X"22",X"03",X"CC",X"00",X"43",X"10",X"83",
		X"00",X"D4",X"25",X"02",X"C6",X"D4",X"34",X"04",X"BD",X"5D",X"BF",X"D6",X"DD",X"58",X"3D",X"1F",
		X"89",X"4F",X"D0",X"DD",X"82",X"00",X"EB",X"35",X"89",X"00",X"2B",X"06",X"10",X"83",X"00",X"11",
		X"22",X"03",X"CC",X"00",X"11",X"10",X"83",X"00",X"7E",X"25",X"02",X"C6",X"7E",X"1F",X"98",X"35",
		X"04",X"84",X"FE",X"C4",X"FC",X"ED",X"4C",X"CC",X"78",X"13",X"ED",X"4A",X"96",X"E3",X"44",X"44",
		X"A7",X"C8",X"16",X"A6",X"5D",X"26",X"07",X"A6",X"5B",X"26",X"03",X"7E",X"74",X"AF",X"10",X"AE",
		X"C8",X"17",X"A6",X"35",X"A0",X"15",X"22",X"01",X"40",X"81",X"19",X"22",X"0E",X"A6",X"37",X"A0",
		X"17",X"22",X"01",X"40",X"81",X"1C",X"22",X"03",X"7E",X"78",X"A9",X"A6",X"C8",X"10",X"A0",X"17",
		X"24",X"01",X"40",X"81",X"04",X"23",X"07",X"86",X"03",X"A7",X"C8",X"11",X"20",X"0F",X"A6",X"C8",
		X"14",X"91",X"D7",X"25",X"2C",X"A6",X"C8",X"11",X"2F",X"27",X"6A",X"C8",X"11",X"A6",X"35",X"A0",
		X"15",X"24",X"01",X"40",X"81",X"01",X"23",X"4C",X"E6",X"37",X"CB",X"05",X"E0",X"17",X"24",X"01",
		X"50",X"54",X"C1",X"01",X"23",X"3E",X"34",X"04",X"A0",X"E0",X"24",X"01",X"40",X"81",X"01",X"23",
		X"33",X"4F",X"E6",X"15",X"C4",X"FE",X"E1",X"4C",X"27",X"08",X"25",X"04",X"8A",X"04",X"20",X"02",
		X"8A",X"08",X"E6",X"17",X"C4",X"FC",X"E1",X"4D",X"27",X"08",X"22",X"04",X"8A",X"02",X"20",X"02",
		X"8A",X"01",X"5F",X"4D",X"27",X"03",X"7E",X"79",X"70",X"6A",X"C8",X"16",X"10",X"2E",X"00",X"AB",
		X"10",X"AE",X"C8",X"17",X"A6",X"35",X"26",X"0A",X"CC",X"00",X"01",X"6D",X"4E",X"27",X"05",X"58",
		X"20",X"02",X"8D",X"18",X"10",X"8E",X"79",X"49",X"10",X"AF",X"4A",X"ED",X"4C",X"96",X"E3",X"A7",
		X"C8",X"16",X"A6",X"17",X"A7",X"C8",X"10",X"A6",X"4C",X"7E",X"79",X"70",X"A6",X"35",X"A0",X"15",
		X"24",X"01",X"40",X"E6",X"37",X"CB",X"05",X"E0",X"17",X"24",X"01",X"50",X"54",X"ED",X"4C",X"A0",
		X"4D",X"24",X"01",X"40",X"A1",X"4C",X"25",X"26",X"E1",X"4C",X"25",X"12",X"E6",X"37",X"CB",X"05",
		X"E1",X"17",X"24",X"05",X"CC",X"40",X"00",X"20",X"3F",X"CC",X"80",X"00",X"20",X"3A",X"E6",X"35",
		X"E1",X"15",X"24",X"05",X"CC",X"00",X"01",X"20",X"2F",X"CC",X"00",X"02",X"20",X"2A",X"A1",X"4D",
		X"22",X"EC",X"E6",X"37",X"CB",X"05",X"E1",X"17",X"25",X"10",X"E6",X"35",X"E1",X"15",X"24",X"05",
		X"CC",X"80",X"01",X"20",X"13",X"CC",X"80",X"02",X"20",X"0E",X"E6",X"35",X"E1",X"15",X"24",X"05",
		X"CC",X"40",X"01",X"20",X"03",X"CC",X"40",X"02",X"39",X"A6",X"5D",X"26",X"13",X"A6",X"5B",X"26",
		X"0F",X"6A",X"C8",X"16",X"2E",X"05",X"CC",X"74",X"AF",X"ED",X"4A",X"4F",X"5F",X"7E",X"79",X"70",
		X"96",X"5C",X"11",X"83",X"99",X"91",X"27",X"02",X"96",X"58",X"84",X"0F",X"E6",X"4D",X"AA",X"4C",
		X"ED",X"C8",X"1A",X"35",X"D0",X"BD",X"D6",X"8B",X"81",X"00",X"00",X"86",X"01",X"BD",X"D6",X"BA",
		X"96",X"22",X"27",X"1E",X"0F",X"39",X"0F",X"68",X"BD",X"D8",X"AB",X"BD",X"D7",X"0D",X"BD",X"7F",
		X"0B",X"CC",X"FF",X"37",X"B7",X"C8",X"0E",X"F7",X"C8",X"0E",X"BD",X"D6",X"8B",X"81",X"BF",X"00",
		X"0F",X"22",X"F6",X"C8",X"04",X"C4",X"30",X"27",X"D2",X"8E",X"CC",X"06",X"BD",X"37",X"BF",X"81",
		X"09",X"27",X"20",X"B6",X"BF",X"32",X"27",X"C3",X"81",X"02",X"24",X"04",X"C5",X"20",X"26",X"BB",
		X"C5",X"20",X"27",X"03",X"8B",X"99",X"19",X"8B",X"99",X"19",X"B7",X"BF",X"32",X"8E",X"CD",X"00",
		X"BD",X"37",X"C8",X"86",X"08",X"0F",X"23",X"C5",X"20",X"27",X"08",X"4C",X"0C",X"23",X"C6",X"0A",
		X"BD",X"37",X"B9",X"1F",X"89",X"BD",X"37",X"B9",X"C6",X"0A",X"BD",X"37",X"B9",X"86",X"02",X"D6",
		X"23",X"27",X"01",X"4F",X"97",X"39",X"CE",X"7A",X"0A",X"AE",X"C1",X"EC",X"C1",X"80",X"6C",X"88",
		X"4A",X"BD",X"46",X"20",X"A6",X"C0",X"26",X"F5",X"20",X"21",X"10",X"F8",X"CC",X"11",X"B3",X"CD",
		X"AC",X"D7",X"C5",X"C8",X"C8",X"C5",X"AD",X"C9",X"C3",X"AC",X"B1",X"C8",X"B1",X"B3",X"C0",X"C2",
		X"BF",X"BE",X"C5",X"B3",X"C3",X"AC",X"C5",X"BE",X"B3",X"D0",X"00",X"BD",X"D7",X"0D",X"BD",X"D8",
		X"5C",X"BD",X"7F",X"0B",X"BD",X"DD",X"0F",X"8E",X"7A",X"9F",X"8D",X"36",X"30",X"04",X"8C",X"7A",
		X"CF",X"25",X"F7",X"CC",X"74",X"11",X"8E",X"30",X"15",X"BD",X"46",X"23",X"10",X"8E",X"7A",X"55",
		X"8D",X"1B",X"7E",X"7B",X"0F",X"75",X"66",X"24",X"30",X"E1",X"99",X"3B",X"65",X"E0",X"22",X"3B",
		X"93",X"E2",X"BB",X"3C",X"C1",X"00",X"E6",X"A0",X"AE",X"A1",X"BD",X"46",X"2C",X"A6",X"A0",X"26",
		X"F5",X"39",X"10",X"AE",X"02",X"A6",X"22",X"E6",X"24",X"E3",X"84",X"10",X"AE",X"A4",X"1A",X"50",
		X"FD",X"CA",X"04",X"EC",X"A4",X"FD",X"CA",X"06",X"31",X"22",X"10",X"BF",X"CA",X"02",X"10",X"AE",
		X"02",X"86",X"0A",X"E6",X"23",X"2A",X"02",X"8A",X"20",X"B7",X"CA",X"00",X"1C",X"AF",X"39",X"45",
		X"56",X"00",X"1C",X"44",X"56",X"07",X"DC",X"45",X"56",X"08",X"FC",X"44",X"56",X"09",X"25",X"45",
		X"84",X"03",X"65",X"44",X"83",X"08",X"24",X"45",X"84",X"09",X"90",X"45",X"84",X"09",X"B9",X"45",
		X"B2",X"04",X"EF",X"44",X"B2",X"08",X"6C",X"45",X"B2",X"09",X"4E",X"45",X"B2",X"09",X"6F",X"45",
		X"B2",X"06",X"41",X"44",X"B2",X"08",X"B4",X"45",X"B2",X"0A",X"28",X"45",X"B2",X"0A",X"49",X"45",
		X"92",X"01",X"D9",X"45",X"92",X"00",X"00",X"45",X"92",X"09",X"E2",X"45",X"92",X"0A",X"05",X"50",
		X"7D",X"AA",X"53",X"80",X"AD",X"34",X"20",X"BD",X"89",X"20",X"A6",X"E0",X"5F",X"ED",X"15",X"ED",
		X"11",X"A6",X"E0",X"ED",X"17",X"A7",X"13",X"EF",X"0A",X"BD",X"D8",X"C6",X"9F",X"2A",X"39",X"DE",
		X"1C",X"CC",X"00",X"50",X"E7",X"4C",X"10",X"8E",X"40",X"4E",X"8D",X"D9",X"AF",X"4D",X"CC",X"00",
		X"FF",X"ED",X"4A",X"96",X"23",X"27",X"0C",X"A7",X"4B",X"86",X"08",X"10",X"8E",X"4C",X"7E",X"8D",
		X"C4",X"AF",X"47",X"86",X"FF",X"97",X"3C",X"0F",X"68",X"96",X"58",X"85",X"30",X"26",X"04",X"0F",
		X"3C",X"20",X"04",X"D6",X"3C",X"27",X"75",X"E6",X"4C",X"C4",X"03",X"10",X"26",X"00",X"62",X"47",
		X"24",X"0D",X"E6",X"4A",X"5A",X"2A",X"02",X"C6",X"02",X"E1",X"4B",X"27",X"F7",X"E7",X"4A",X"47",
		X"24",X"0E",X"E6",X"4A",X"5C",X"C1",X"03",X"26",X"01",X"5F",X"E1",X"4B",X"27",X"F6",X"E7",X"4A",
		X"D6",X"5C",X"57",X"24",X"0F",X"A6",X"4B",X"2B",X"1E",X"4A",X"2A",X"02",X"86",X"02",X"A1",X"4A",
		X"27",X"F7",X"A7",X"4B",X"57",X"24",X"10",X"A6",X"4B",X"2B",X"0C",X"4C",X"81",X"03",X"26",X"01",
		X"4F",X"A1",X"4A",X"27",X"F6",X"A7",X"4B",X"A6",X"4A",X"10",X"8E",X"7A",X"EF",X"A6",X"A6",X"AE",
		X"4D",X"A7",X"17",X"A6",X"4B",X"2B",X"0A",X"10",X"8E",X"7A",X"F2",X"A6",X"A6",X"AE",X"47",X"A7",
		X"17",X"86",X"05",X"BD",X"D6",X"BA",X"6A",X"4C",X"10",X"26",X"FF",X"7B",X"BD",X"D8",X"AB",X"BD",
		X"7F",X"0B",X"1A",X"F0",X"DE",X"1C",X"A6",X"4A",X"CE",X"99",X"91",X"C6",X"01",X"8E",X"25",X"48",
		X"BD",X"7C",X"60",X"DE",X"1C",X"A6",X"4B",X"2A",X"02",X"86",X"03",X"CE",X"99",X"D9",X"C6",X"02",
		X"8E",X"70",X"48",X"BD",X"7C",X"60",X"96",X"23",X"26",X"14",X"BE",X"99",X"CC",X"A7",X"11",X"BE",
		X"99",X"CE",X"A7",X"11",X"BE",X"99",X"D2",X"A7",X"11",X"BE",X"99",X"D0",X"A7",X"11",X"BD",X"D6",
		X"8B",X"E9",X"D6",X"28",X"CE",X"9A",X"21",X"4F",X"5F",X"ED",X"C8",X"27",X"4C",X"ED",X"53",X"10",
		X"8E",X"7A",X"DF",X"86",X"04",X"A7",X"C8",X"25",X"8D",X"34",X"34",X"20",X"10",X"8E",X"25",X"88",
		X"BD",X"D8",X"8E",X"6F",X"11",X"AF",X"55",X"35",X"20",X"31",X"24",X"8D",X"21",X"CC",X"25",X"88",
		X"BD",X"7C",X"E0",X"86",X"80",X"A7",X"19",X"6F",X"11",X"AF",X"57",X"8D",X"11",X"CC",X"25",X"88",
		X"BD",X"7C",X"E0",X"86",X"81",X"A7",X"19",X"6F",X"11",X"AF",X"59",X"7E",X"7D",X"24",X"BD",X"D7",
		X"50",X"6C",X"02",X"EF",X"0A",X"EC",X"22",X"ED",X"08",X"86",X"08",X"A7",X"03",X"31",X"24",X"39",
		X"34",X"34",X"A7",X"C8",X"25",X"C6",X"10",X"3D",X"10",X"8E",X"7A",X"9F",X"31",X"A5",X"86",X"44",
		X"E6",X"E4",X"56",X"25",X"02",X"86",X"22",X"34",X"02",X"BD",X"7D",X"00",X"10",X"AF",X"64",X"10",
		X"AE",X"62",X"BD",X"D8",X"8E",X"AF",X"55",X"10",X"AE",X"64",X"BD",X"7D",X"00",X"10",X"AF",X"64",
		X"EC",X"62",X"8D",X"4C",X"86",X"C0",X"A7",X"19",X"AF",X"53",X"BD",X"7D",X"00",X"10",X"AF",X"64",
		X"EC",X"62",X"8D",X"3C",X"86",X"80",X"A7",X"19",X"AF",X"57",X"10",X"AE",X"64",X"BD",X"7D",X"00",
		X"EC",X"62",X"8D",X"2C",X"86",X"81",X"A7",X"19",X"AF",X"59",X"35",X"B6",X"34",X"24",X"20",X"10",
		X"34",X"24",X"5F",X"10",X"AE",X"08",X"E3",X"22",X"ED",X"11",X"ED",X"15",X"A6",X"E4",X"AB",X"24",
		X"A7",X"13",X"5F",X"ED",X"17",X"E7",X"04",X"E7",X"05",X"E7",X"02",X"BD",X"D8",X"C6",X"35",X"A4",
		X"34",X"24",X"5F",X"10",X"AE",X"08",X"E3",X"22",X"ED",X"11",X"ED",X"15",X"A6",X"E4",X"AB",X"24",
		X"A7",X"13",X"5F",X"ED",X"17",X"E7",X"04",X"E7",X"05",X"BD",X"D8",X"C6",X"9F",X"2A",X"35",X"A4",
		X"BD",X"D7",X"50",X"EF",X"0A",X"EC",X"22",X"ED",X"08",X"EC",X"62",X"A7",X"0C",X"E7",X"03",X"31",
		X"24",X"39",X"67",X"44",X"25",X"0F",X"DF",X"22",X"32",X"0D",X"00",X"67",X"44",X"65",X"0F",X"DF",
		X"22",X"58",X"0D",X"00",X"1C",X"AF",X"BD",X"DD",X"0F",X"CC",X"5E",X"DD",X"8E",X"06",X"13",X"BD",
		X"46",X"23",X"10",X"8E",X"7D",X"12",X"BD",X"7A",X"6D",X"96",X"23",X"27",X"0C",X"CC",X"5F",X"DD",
		X"8E",X"78",X"13",X"BD",X"46",X"23",X"BD",X"7A",X"6D",X"4F",X"5F",X"FD",X"99",X"BC",X"FD",X"99",
		X"BE",X"FD",X"9A",X"04",X"FD",X"9A",X"06",X"FD",X"9A",X"4C",X"FD",X"9A",X"4E",X"1A",X"50",X"CC",
		X"90",X"1B",X"FD",X"CA",X"04",X"86",X"FF",X"B7",X"CA",X"01",X"C6",X"CC",X"86",X"07",X"FD",X"CA",
		X"06",X"C6",X"32",X"F7",X"CA",X"00",X"8E",X"00",X"1B",X"BF",X"CA",X"04",X"C6",X"FF",X"F7",X"CA",
		X"01",X"86",X"06",X"C6",X"CD",X"FD",X"CA",X"06",X"C6",X"12",X"F7",X"CA",X"00",X"8E",X"05",X"1B",
		X"BF",X"CA",X"04",X"86",X"FF",X"B7",X"CA",X"01",X"C6",X"01",X"86",X"8C",X"FD",X"CA",X"06",X"C6",
		X"12",X"F7",X"CA",X"00",X"86",X"95",X"C6",X"18",X"FD",X"CA",X"06",X"8E",X"00",X"E7",X"BF",X"CA",
		X"04",X"C6",X"12",X"F7",X"CA",X"00",X"8E",X"CC",X"14",X"BD",X"37",X"BF",X"6F",X"E2",X"81",X"03",
		X"23",X"08",X"6C",X"E4",X"81",X"06",X"23",X"02",X"6C",X"E4",X"8E",X"64",X"DE",X"10",X"8E",X"98",
		X"D3",X"E6",X"E4",X"58",X"EC",X"85",X"ED",X"A4",X"86",X"02",X"A7",X"22",X"30",X"0E",X"31",X"23",
		X"8C",X"65",X"E8",X"25",X"EC",X"32",X"61",X"B6",X"99",X"04",X"97",X"D0",X"CC",X"02",X"00",X"FD",
		X"99",X"96",X"FD",X"99",X"DE",X"FD",X"9A",X"26",X"CC",X"01",X"00",X"FD",X"99",X"94",X"FD",X"99",
		X"DC",X"FD",X"9A",X"24",X"8E",X"CC",X"02",X"BD",X"37",X"BF",X"B7",X"99",X"11",X"B7",X"99",X"1A",
		X"8E",X"CC",X"04",X"BD",X"37",X"C2",X"4F",X"58",X"49",X"58",X"49",X"58",X"49",X"58",X"49",X"DD",
		X"B8",X"FD",X"99",X"13",X"FD",X"99",X"1C",X"8E",X"CC",X"00",X"BD",X"37",X"C2",X"BD",X"37",X"DD",
		X"86",X"87",X"3D",X"58",X"49",X"97",X"8B",X"97",X"8C",X"4F",X"BD",X"E7",X"FD",X"97",X"73",X"97",
		X"87",X"B7",X"BF",X"34",X"B6",X"99",X"07",X"97",X"BB",X"97",X"85",X"86",X"2C",X"97",X"BA",X"CC",
		X"07",X"07",X"DD",X"CC",X"CC",X"6A",X"B3",X"DD",X"CE",X"CE",X"99",X"91",X"BD",X"74",X"15",X"CE",
		X"99",X"D9",X"BD",X"74",X"15",X"CE",X"9A",X"21",X"BD",X"74",X"15",X"86",X"80",X"9A",X"39",X"97",
		X"39",X"48",X"2B",X"06",X"BD",X"D6",X"8B",X"5F",X"8D",X"56",X"BD",X"D6",X"8B",X"E2",X"3A",X"10",
		X"BD",X"D6",X"8B",X"E5",X"46",X"12",X"BD",X"D6",X"8B",X"E7",X"9A",X"15",X"BD",X"D6",X"8B",X"DD",
		X"3F",X"14",X"86",X"04",X"97",X"8E",X"86",X"40",X"97",X"8F",X"BD",X"D6",X"8B",X"E7",X"13",X"13",
		X"6C",X"04",X"BD",X"D6",X"8B",X"65",X"E8",X"16",X"6C",X"04",X"CC",X"68",X"2F",X"ED",X"07",X"86",
		X"1F",X"8B",X"14",X"A7",X"09",X"8B",X"14",X"A7",X"0B",X"BD",X"5D",X"BF",X"84",X"3F",X"8B",X"28",
		X"A7",X"0C",X"86",X"FF",X"A7",X"0A",X"96",X"23",X"27",X"0A",X"97",X"86",X"BD",X"D6",X"8B",X"E2",
		X"41",X"11",X"6C",X"04",X"BD",X"D6",X"8B",X"E9",X"89",X"20",X"6C",X"04",X"6C",X"04",X"BD",X"D6",
		X"8B",X"60",X"00",X"17",X"6C",X"04",X"6C",X"04",X"CC",X"1B",X"DB",X"ED",X"09",X"CE",X"98",X"90",
		X"EF",X"0D",X"BD",X"D6",X"8B",X"60",X"00",X"18",X"A6",X"04",X"8B",X"03",X"A7",X"04",X"86",X"6C",
		X"ED",X"09",X"33",X"41",X"EF",X"0D",X"1C",X"AF",X"7E",X"D6",X"C5",X"1A",X"50",X"BD",X"D8",X"6D",
		X"BD",X"D8",X"F1",X"1C",X"AF",X"BD",X"DD",X"0F",X"7E",X"D8",X"5C",X"0F",X"39",X"96",X"39",X"26",
		X"0E",X"BD",X"D8",X"AB",X"BD",X"D7",X"0D",X"8D",X"E2",X"BD",X"D6",X"8B",X"79",X"75",X"00",X"7E",
		X"D6",X"C5",X"0F",X"39",X"8D",X"D5",X"86",X"4A",X"97",X"05",X"86",X"03",X"BD",X"D6",X"BA",X"BD",
		X"DE",X"44",X"CC",X"5B",X"88",X"8E",X"1A",X"C0",X"BD",X"46",X"23",X"BD",X"37",X"E3",X"BD",X"E3",
		X"52",X"DE",X"1C",X"86",X"03",X"A7",X"47",X"86",X"A0",X"BD",X"D6",X"BA",X"6A",X"47",X"26",X"F7",
		X"BD",X"D8",X"AB",X"BD",X"D7",X"0D",X"8D",X"A3",X"BD",X"D6",X"8B",X"80",X"ED",X"50",X"BD",X"D6",
		X"8B",X"79",X"7B",X"24",X"DE",X"1C",X"10",X"8E",X"80",X"16",X"10",X"AF",X"48",X"86",X"1E",X"BD",
		X"D6",X"BA",X"86",X"60",X"97",X"8B",X"4F",X"5F",X"DD",X"B8",X"10",X"AE",X"48",X"EC",X"A1",X"10",
		X"2B",X"FF",X"88",X"10",X"AF",X"48",X"E7",X"47",X"8E",X"7F",X"BD",X"AD",X"86",X"10",X"AE",X"48",
		X"BD",X"7A",X"6D",X"86",X"04",X"BD",X"D6",X"BA",X"6A",X"47",X"26",X"F1",X"10",X"AE",X"48",X"A6",
		X"A0",X"27",X"C7",X"31",X"21",X"5F",X"AE",X"A1",X"BD",X"46",X"2C",X"20",X"F2",X"03",X"73",X"86",
		X"01",X"97",X"83",X"0F",X"85",X"0C",X"86",X"8E",X"80",X"06",X"86",X"26",X"BD",X"D6",X"76",X"20",
		X"0C",X"86",X"25",X"8E",X"82",X"C8",X"BD",X"D6",X"76",X"0C",X"74",X"0C",X"88",X"BD",X"D6",X"8B",
		X"81",X"E5",X"23",X"86",X"04",X"A7",X"08",X"39",X"0F",X"83",X"0F",X"86",X"8E",X"60",X"CE",X"86",
		X"29",X"BD",X"D6",X"76",X"CC",X"1D",X"E7",X"ED",X"07",X"0F",X"D1",X"39",X"0C",X"D1",X"0C",X"85",
		X"39",X"86",X"05",X"97",X"73",X"39",X"8E",X"86",X"1C",X"86",X"26",X"BD",X"D6",X"76",X"86",X"78",
		X"BD",X"D6",X"BA",X"7E",X"86",X"1C",X"3E",X"5A",X"FF",X"33",X"2C",X"C0",X"FE",X"22",X"2C",X"C8",
		X"FD",X"22",X"2C",X"D0",X"00",X"3E",X"4B",X"FC",X"22",X"20",X"C8",X"FB",X"22",X"20",X"D0",X"00",
		X"3E",X"4B",X"FA",X"22",X"22",X"C8",X"F9",X"22",X"22",X"D0",X"00",X"3E",X"69",X"C9",X"22",X"22",
		X"C8",X"CA",X"22",X"26",X"D0",X"CB",X"22",X"22",X"D8",X"CC",X"22",X"26",X"E0",X"00",X"14",X"4B",
		X"F8",X"22",X"26",X"C8",X"F7",X"22",X"26",X"D0",X"00",X"44",X"4B",X"E9",X"22",X"23",X"C8",X"E8",
		X"22",X"23",X"D0",X"00",X"00",X"69",X"E7",X"22",X"2C",X"C8",X"DE",X"22",X"2F",X"D0",X"DD",X"22",
		X"2C",X"D8",X"DC",X"22",X"2F",X"E0",X"00",X"2B",X"69",X"D7",X"22",X"2B",X"C8",X"04",X"22",X"2F",
		X"D0",X"03",X"22",X"2B",X"D8",X"02",X"22",X"2F",X"E0",X"00",X"3F",X"69",X"DB",X"22",X"26",X"C8",
		X"DA",X"22",X"2A",X"D0",X"D9",X"22",X"26",X"D8",X"D8",X"22",X"2A",X"E0",X"00",X"3E",X"5A",X"F6",
		X"11",X"2B",X"98",X"F5",X"44",X"2B",X"A0",X"F3",X"44",X"2B",X"A8",X"F4",X"44",X"2B",X"B0",X"F2",
		X"44",X"2B",X"B8",X"F1",X"44",X"2B",X"C0",X"F0",X"44",X"2B",X"C8",X"01",X"44",X"2B",X"D0",X"E5",
		X"44",X"2B",X"D8",X"E4",X"22",X"2B",X"E0",X"EF",X"44",X"66",X"A0",X"EE",X"44",X"66",X"A8",X"ED",
		X"44",X"66",X"B0",X"EC",X"44",X"66",X"B8",X"ED",X"44",X"66",X"C0",X"EA",X"44",X"66",X"C8",X"EB",
		X"44",X"66",X"D0",X"EB",X"44",X"66",X"D8",X"E6",X"22",X"66",X"E0",X"00",X"FF",X"1A",X"50",X"86",
		X"42",X"97",X"39",X"0F",X"23",X"4F",X"5F",X"FD",X"99",X"82",X"5C",X"ED",X"4A",X"7E",X"7B",X"C4",
		X"0F",X"68",X"0F",X"39",X"BD",X"7F",X"0B",X"86",X"03",X"BD",X"D6",X"BA",X"86",X"0F",X"A7",X"47",
		X"BD",X"37",X"D1",X"BD",X"D6",X"8B",X"81",X"3A",X"00",X"86",X"32",X"BD",X"D6",X"BA",X"6A",X"47",
		X"26",X"F1",X"86",X"03",X"ED",X"47",X"86",X"FE",X"BD",X"D6",X"BA",X"6A",X"47",X"26",X"F7",X"8E",
		X"7F",X"32",X"A6",X"45",X"BD",X"D6",X"76",X"7E",X"D6",X"C5",X"BD",X"5D",X"BF",X"C6",X"05",X"3D",
		X"48",X"BD",X"D7",X"50",X"A7",X"19",X"48",X"10",X"8E",X"00",X"00",X"10",X"AE",X"A6",X"10",X"AF",
		X"08",X"10",X"AE",X"A4",X"31",X"22",X"10",X"AF",X"1A",X"C6",X"D0",X"EB",X"3E",X"E7",X"14",X"86",
		X"04",X"A7",X"03",X"CC",X"86",X"00",X"ED",X"15",X"ED",X"11",X"86",X"D0",X"ED",X"17",X"A7",X"13",
		X"4F",X"ED",X"1C",X"CC",X"FE",X"FF",X"ED",X"1E",X"AF",X"47",X"EF",X"0A",X"9F",X"2A",X"86",X"01",
		X"BD",X"D6",X"BA",X"AE",X"47",X"A6",X"11",X"26",X"06",X"BD",X"D7",X"84",X"7E",X"D6",X"C5",X"86",
		X"DA",X"A1",X"17",X"22",X"0A",X"4F",X"5F",X"ED",X"1E",X"C6",X"80",X"ED",X"1C",X"20",X"DF",X"86",
		X"08",X"A1",X"15",X"25",X"09",X"4F",X"5F",X"ED",X"1C",X"4C",X"ED",X"1E",X"20",X"D0",X"86",X"54",
		X"A1",X"17",X"25",X"CA",X"4F",X"5F",X"ED",X"1E",X"CC",X"FF",X"80",X"ED",X"1C",X"20",X"BF",X"86",
		X"30",X"A7",X"49",X"86",X"12",X"F6",X"BF",X"32",X"5A",X"27",X"02",X"86",X"13",X"BD",X"46",X"32",
		X"BD",X"E3",X"52",X"86",X"F4",X"BD",X"D6",X"BA",X"6A",X"49",X"26",X"F7",X"BD",X"D6",X"8B",X"81",
		X"00",X"00",X"7E",X"D6",X"C5",X"8E",X"98",X"01",X"C6",X"FF",X"E7",X"80",X"8C",X"98",X"10",X"26",
		X"F9",X"C6",X"04",X"E7",X"47",X"86",X"05",X"BD",X"D6",X"BA",X"BD",X"D8",X"5C",X"86",X"1E",X"BD",
		X"D6",X"BA",X"A6",X"48",X"BD",X"E9",X"72",X"86",X"05",X"BD",X"D6",X"BA",X"86",X"08",X"BD",X"89",
		X"20",X"A6",X"48",X"48",X"48",X"10",X"8E",X"82",X"9C",X"31",X"A6",X"A6",X"A0",X"5F",X"ED",X"15",
		X"ED",X"11",X"A6",X"A0",X"ED",X"17",X"A7",X"13",X"CC",X"01",X"2F",X"8D",X"34",X"47",X"56",X"ED",
		X"1C",X"CC",X"01",X"2F",X"8D",X"2B",X"ED",X"1E",X"BD",X"D8",X"C6",X"31",X"84",X"BD",X"D6",X"8B",
		X"6C",X"01",X"22",X"10",X"AF",X"07",X"AF",X"2A",X"10",X"9F",X"2A",X"6A",X"47",X"27",X"08",X"86",
		X"06",X"8E",X"82",X"0C",X"7E",X"D6",X"BC",X"A6",X"48",X"8E",X"98",X"A3",X"6A",X"86",X"7E",X"D6",
		X"C5",X"A7",X"E2",X"BD",X"5D",X"BF",X"A7",X"E2",X"3D",X"AB",X"61",X"6D",X"A0",X"2E",X"0A",X"2D",
		X"04",X"64",X"E4",X"24",X"04",X"43",X"50",X"82",X"FF",X"32",X"62",X"47",X"56",X"47",X"56",X"47",
		X"56",X"47",X"56",X"39",X"10",X"8E",X"82",X"B2",X"CC",X"10",X"20",X"8D",X"D4",X"47",X"56",X"ED",
		X"1C",X"CC",X"10",X"20",X"BD",X"82",X"61",X"ED",X"1E",X"7E",X"D8",X"C6",X"07",X"BB",X"01",X"00",
		X"07",X"50",X"01",X"00",X"88",X"50",X"FF",X"00",X"88",X"BB",X"FF",X"00",X"49",X"39",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"02",X"80",X"03",X"01",X"01",X"00",X"02",
		X"02",X"01",X"80",X"03",X"01",X"01",X"00",X"02",X"86",X"04",X"BD",X"E9",X"72",X"86",X"05",X"BD",
		X"D6",X"BA",X"CC",X"0A",X"0F",X"A7",X"C8",X"35",X"E7",X"C8",X"37",X"CC",X"82",X"E7",X"ED",X"C8",
		X"38",X"CC",X"1F",X"42",X"7E",X"85",X"A6",X"BD",X"D7",X"3C",X"1E",X"A0",X"00",X"9F",X"7E",X"86",
		X"40",X"A7",X"03",X"AF",X"47",X"CC",X"44",X"00",X"ED",X"15",X"CC",X"39",X"00",X"ED",X"17",X"CC",
		X"44",X"00",X"ED",X"11",X"86",X"35",X"A7",X"13",X"BD",X"D8",X"C6",X"86",X"10",X"A7",X"19",X"9F",
		X"2A",X"6F",X"4A",X"0A",X"88",X"96",X"75",X"10",X"26",X"01",X"6B",X"86",X"01",X"03",X"80",X"2A",
		X"01",X"40",X"A7",X"4D",X"6F",X"49",X"86",X"07",X"A7",X"4E",X"BD",X"84",X"37",X"A6",X"4E",X"8E",
		X"83",X"35",X"7E",X"D6",X"BC",X"BD",X"84",X"4A",X"DE",X"1C",X"BD",X"8A",X"DC",X"48",X"48",X"10",
		X"8E",X"82",X"B8",X"31",X"A6",X"EC",X"21",X"6D",X"4D",X"2A",X"04",X"43",X"50",X"82",X"FF",X"E3",
		X"15",X"81",X"1D",X"24",X"04",X"86",X"1D",X"20",X"5D",X"81",X"6F",X"25",X"04",X"86",X"6F",X"20",
		X"55",X"ED",X"15",X"A6",X"23",X"AB",X"17",X"81",X"D6",X"24",X"04",X"A7",X"17",X"20",X"BB",X"86",
		X"FF",X"A7",X"03",X"86",X"02",X"BD",X"D6",X"BA",X"AE",X"47",X"6C",X"02",X"A6",X"11",X"27",X"03",
		X"BD",X"DC",X"73",X"31",X"84",X"0F",X"7E",X"0F",X"7F",X"BD",X"D6",X"8B",X"89",X"7A",X"00",X"A6",
		X"35",X"C6",X"DA",X"ED",X"07",X"CC",X"1F",X"6E",X"ED",X"09",X"FC",X"1F",X"6C",X"ED",X"0B",X"6F",
		X"0D",X"86",X"05",X"A7",X"0E",X"86",X"14",X"BD",X"D6",X"BA",X"0A",X"74",X"AE",X"47",X"BD",X"D7",
		X"84",X"0F",X"C9",X"7E",X"D6",X"C5",X"A7",X"15",X"86",X"01",X"A7",X"05",X"BD",X"84",X"4A",X"27",
		X"09",X"8D",X"1F",X"86",X"0A",X"BD",X"D6",X"BA",X"8D",X"36",X"DE",X"1C",X"BD",X"84",X"37",X"4D",
		X"10",X"26",X"FF",X"56",X"96",X"C9",X"27",X"02",X"6C",X"0C",X"86",X"02",X"8E",X"83",X"BC",X"7E",
		X"D6",X"BC",X"DE",X"1C",X"AE",X"47",X"86",X"03",X"A7",X"05",X"86",X"05",X"AB",X"17",X"A7",X"17",
		X"AE",X"06",X"A6",X"19",X"84",X"0E",X"A7",X"C8",X"1B",X"8E",X"E6",X"64",X"BD",X"E6",X"AA",X"39",
		X"AE",X"47",X"86",X"01",X"A7",X"05",X"A6",X"17",X"80",X"05",X"A7",X"17",X"81",X"3F",X"25",X"26",
		X"A6",X"15",X"8B",X"02",X"E6",X"17",X"C0",X"06",X"DD",X"43",X"10",X"8E",X"82",X"B6",X"CC",X"08",
		X"00",X"BD",X"82",X"61",X"DD",X"3F",X"CC",X"10",X"10",X"BD",X"82",X"61",X"DD",X"41",X"A6",X"C8",
		X"1B",X"C6",X"C4",X"BD",X"88",X"E4",X"39",X"AE",X"47",X"A6",X"0C",X"27",X"0A",X"E6",X"49",X"26",
		X"08",X"60",X"4D",X"86",X"02",X"A7",X"4E",X"A7",X"49",X"39",X"AE",X"47",X"10",X"AE",X"1A",X"EC",
		X"11",X"10",X"83",X"25",X"00",X"25",X"07",X"CC",X"70",X"00",X"A0",X"3E",X"20",X"13",X"CC",X"1E",
		X"00",X"A0",X"3E",X"10",X"A3",X"11",X"22",X"06",X"33",X"84",X"BD",X"D2",X"B1",X"39",X"C3",X"52",
		X"00",X"10",X"A3",X"11",X"22",X"0E",X"CC",X"77",X"00",X"10",X"A3",X"11",X"23",X"06",X"33",X"84",
		X"BD",X"D2",X"D2",X"39",X"5F",X"39",X"6F",X"03",X"CC",X"85",X"44",X"ED",X"4B",X"86",X"0A",X"A7",
		X"C8",X"11",X"CC",X"83",X"A5",X"ED",X"4D",X"CC",X"84",X"D2",X"ED",X"C8",X"13",X"CC",X"85",X"89",
		X"ED",X"C8",X"15",X"C6",X"02",X"8D",X"60",X"7E",X"85",X"DF",X"86",X"05",X"A7",X"C8",X"17",X"96",
		X"75",X"26",X"16",X"C1",X"D5",X"10",X"24",X"FE",X"B6",X"CC",X"86",X"0E",X"ED",X"C8",X"13",X"86",
		X"03",X"A7",X"C8",X"11",X"CC",X"00",X"06",X"20",X"DE",X"86",X"07",X"A7",X"C8",X"11",X"8D",X"08",
		X"20",X"D5",X"6F",X"0C",X"86",X"01",X"20",X"F3",X"10",X"8E",X"98",X"3F",X"A6",X"15",X"80",X"06",
		X"A7",X"A0",X"86",X"9A",X"A0",X"15",X"A7",X"A0",X"A6",X"17",X"80",X"37",X"47",X"A7",X"A0",X"86",
		X"F6",X"A0",X"17",X"47",X"A7",X"A0",X"C6",X"03",X"86",X"FF",X"A1",X"A2",X"25",X"04",X"A6",X"A4",
		X"D7",X"3C",X"5A",X"2A",X"F5",X"D6",X"3C",X"86",X"0A",X"3D",X"D7",X"3C",X"BD",X"5D",X"BF",X"C6",
		X"05",X"3D",X"48",X"9B",X"3C",X"10",X"8E",X"85",X"1C",X"EC",X"A6",X"39",X"01",X"FC",X"02",X"FE",
		X"03",X"00",X"02",X"02",X"01",X"04",X"FF",X"FC",X"FE",X"FE",X"FD",X"00",X"FE",X"02",X"FF",X"04",
		X"FE",X"02",X"FF",X"04",X"00",X"06",X"01",X"04",X"02",X"02",X"FE",X"FE",X"FF",X"FC",X"00",X"FA",
		X"01",X"FC",X"02",X"FE",X"BD",X"8A",X"DC",X"6A",X"C8",X"17",X"26",X"2F",X"A6",X"06",X"27",X"1C",
		X"10",X"AE",X"06",X"A6",X"39",X"81",X"10",X"26",X"13",X"10",X"AC",X"C8",X"1E",X"27",X"09",X"60",
		X"4F",X"60",X"C8",X"10",X"10",X"AF",X"C8",X"1E",X"6F",X"06",X"20",X"03",X"6F",X"C8",X"1E",X"BD",
		X"84",X"4A",X"26",X"08",X"DE",X"1C",X"AE",X"47",X"6C",X"C8",X"17",X"39",X"BD",X"83",X"E2",X"86",
		X"0A",X"BD",X"D6",X"BA",X"BD",X"84",X"00",X"20",X"60",X"A6",X"15",X"E6",X"17",X"81",X"0C",X"10",
		X"25",X"FF",X"17",X"81",X"7B",X"10",X"24",X"FF",X"11",X"C1",X"43",X"10",X"25",X"FF",X"0B",X"C1",
		X"CD",X"10",X"24",X"FF",X"05",X"39",X"6F",X"C8",X"34",X"6F",X"C8",X"36",X"ED",X"C8",X"3A",X"1A",
		X"50",X"FD",X"CA",X"02",X"CC",X"44",X"35",X"FD",X"CA",X"04",X"6C",X"C8",X"36",X"EC",X"C8",X"35",
		X"FD",X"CA",X"06",X"86",X"02",X"B7",X"CA",X"00",X"1C",X"AF",X"E1",X"C8",X"37",X"27",X"0D",X"86",
		X"01",X"BD",X"D6",X"BA",X"EC",X"C8",X"3A",X"A3",X"C8",X"34",X"20",X"D0",X"6E",X"D8",X"38",X"ED",
		X"4F",X"A6",X"C8",X"11",X"A7",X"C8",X"12",X"6F",X"02",X"AE",X"47",X"A6",X"0C",X"26",X"27",X"A6",
		X"11",X"27",X"26",X"6A",X"C8",X"12",X"26",X"16",X"A6",X"C8",X"11",X"A7",X"C8",X"12",X"AD",X"D8",
		X"0B",X"EC",X"4F",X"AB",X"15",X"EB",X"17",X"A7",X"15",X"E7",X"17",X"AD",X"D8",X"15",X"86",X"01",
		X"8E",X"85",X"E9",X"7E",X"D6",X"BC",X"6E",X"D8",X"13",X"6E",X"D8",X"0D",X"6F",X"4A",X"BD",X"EA",
		X"FA",X"2A",X"02",X"86",X"04",X"A7",X"4C",X"BD",X"E9",X"72",X"81",X"04",X"27",X"0F",X"86",X"03",
		X"A0",X"4C",X"BD",X"E9",X"72",X"86",X"14",X"8E",X"86",X"57",X"7E",X"D6",X"BC",X"86",X"05",X"BD",
		X"D6",X"BA",X"CC",X"09",X"13",X"A7",X"C8",X"35",X"E7",X"C8",X"37",X"CC",X"86",X"57",X"ED",X"C8",
		X"38",X"CC",X"21",X"FD",X"7E",X"85",X"A6",X"BD",X"D7",X"3C",X"21",X"4A",X"00",X"AF",X"47",X"A6",
		X"4C",X"48",X"10",X"8E",X"89",X"70",X"31",X"A6",X"81",X"08",X"A6",X"21",X"A7",X"13",X"25",X"02",
		X"8B",X"02",X"ED",X"17",X"A6",X"A4",X"5F",X"ED",X"11",X"ED",X"15",X"C6",X"84",X"E7",X"03",X"BD",
		X"D8",X"C6",X"86",X"20",X"A7",X"19",X"9F",X"2A",X"E6",X"4C",X"CE",X"03",X"80",X"C1",X"04",X"26",
		X"06",X"EF",X"1E",X"86",X"01",X"20",X"11",X"CE",X"FD",X"00",X"C1",X"01",X"23",X"04",X"86",X"02",
		X"20",X"04",X"CE",X"03",X"00",X"4F",X"EF",X"1C",X"A7",X"05",X"8E",X"E6",X"7B",X"BD",X"E6",X"AA",
		X"BD",X"5D",X"BF",X"C6",X"17",X"3D",X"8A",X"04",X"8E",X"86",X"BE",X"7E",X"D6",X"BC",X"AE",X"47",
		X"4F",X"5F",X"ED",X"1C",X"ED",X"1E",X"1A",X"50",X"A6",X"11",X"BD",X"88",X"BE",X"A7",X"15",X"A6",
		X"13",X"BD",X"88",X"D1",X"A7",X"17",X"1C",X"AF",X"A6",X"11",X"10",X"27",X"01",X"8B",X"A6",X"0C",
		X"10",X"26",X"01",X"32",X"96",X"F8",X"A7",X"4B",X"BE",X"99",X"86",X"03",X"7C",X"2A",X"03",X"BE",
		X"99",X"CE",X"AF",X"4D",X"6F",X"4C",X"6F",X"C8",X"11",X"86",X"02",X"BD",X"D6",X"BA",X"6F",X"4F",
		X"6F",X"C8",X"10",X"AE",X"4D",X"10",X"AE",X"47",X"A6",X"2C",X"10",X"26",X"01",X"08",X"A6",X"35",
		X"E6",X"33",X"DD",X"BD",X"BD",X"89",X"35",X"91",X"FB",X"25",X"04",X"6F",X"4C",X"20",X"34",X"91",
		X"FE",X"24",X"04",X"6C",X"4F",X"20",X"2C",X"EC",X"15",X"A3",X"35",X"2A",X"04",X"43",X"50",X"82",
		X"FF",X"48",X"48",X"97",X"3C",X"EC",X"17",X"A3",X"37",X"2A",X"04",X"43",X"50",X"82",X"FF",X"91",
		X"3C",X"24",X"76",X"A6",X"4C",X"26",X"0C",X"A6",X"37",X"81",X"85",X"25",X"04",X"86",X"7F",X"A7",
		X"4C",X"6C",X"4C",X"AE",X"47",X"10",X"AE",X"4D",X"CE",X"99",X"91",X"10",X"BC",X"99",X"86",X"27",
		X"03",X"CE",X"99",X"D9",X"BD",X"6B",X"F3",X"DE",X"1C",X"10",X"25",X"00",X"63",X"A6",X"15",X"E6",
		X"31",X"10",X"27",X"00",X"5B",X"A1",X"31",X"E6",X"4F",X"27",X"04",X"25",X"06",X"20",X"02",X"24",
		X"02",X"8B",X"04",X"80",X"02",X"BD",X"88",X"BE",X"A7",X"15",X"E6",X"17",X"6D",X"4C",X"27",X"04",
		X"2A",X"0E",X"20",X"0E",X"E1",X"33",X"A6",X"4F",X"27",X"04",X"25",X"06",X"20",X"02",X"24",X"02",
		X"CB",X"06",X"C0",X"03",X"BD",X"88",X"D1",X"E7",X"17",X"BD",X"89",X"5D",X"A6",X"4F",X"10",X"27",
		X"FF",X"47",X"A6",X"C8",X"10",X"10",X"27",X"FF",X"40",X"CC",X"06",X"84",X"DD",X"45",X"10",X"AE",
		X"4D",X"A6",X"35",X"E6",X"37",X"C0",X"08",X"DD",X"47",X"BD",X"88",X"78",X"6A",X"4B",X"26",X"1A",
		X"A6",X"C8",X"11",X"26",X"1B",X"6C",X"C8",X"11",X"96",X"F8",X"A7",X"4B",X"FC",X"99",X"CE",X"10",
		X"BC",X"99",X"86",X"27",X"03",X"FC",X"99",X"86",X"ED",X"4D",X"B6",X"99",X"01",X"7E",X"86",X"FB",
		X"AE",X"47",X"86",X"FF",X"E6",X"11",X"C1",X"45",X"24",X"02",X"86",X"01",X"A7",X"49",X"A6",X"15",
		X"AB",X"49",X"A7",X"15",X"BD",X"89",X"5D",X"86",X"01",X"BD",X"D6",X"BA",X"AE",X"47",X"A6",X"11",
		X"27",X"04",X"A6",X"0C",X"27",X"E8",X"AE",X"47",X"A6",X"11",X"26",X"09",X"A6",X"15",X"BD",X"88",
		X"BE",X"A7",X"15",X"A7",X"11",X"86",X"FF",X"A7",X"03",X"86",X"02",X"BD",X"D6",X"BA",X"AE",X"47",
		X"6C",X"02",X"BD",X"DC",X"73",X"31",X"84",X"BD",X"D6",X"8B",X"89",X"7A",X"21",X"A6",X"35",X"E6",
		X"37",X"BD",X"88",X"BE",X"BD",X"88",X"D1",X"ED",X"07",X"CC",X"22",X"30",X"ED",X"09",X"FC",X"22",
		X"2E",X"ED",X"0B",X"33",X"84",X"86",X"FF",X"E6",X"2C",X"27",X"0A",X"0C",X"7D",X"8E",X"E6",X"86",
		X"BD",X"E6",X"AA",X"86",X"44",X"C6",X"05",X"ED",X"4D",X"86",X"14",X"BD",X"D6",X"BA",X"AE",X"47",
		X"0A",X"7B",X"BD",X"D7",X"84",X"7E",X"D6",X"C5",X"AE",X"47",X"A6",X"15",X"E6",X"17",X"CB",X"06",
		X"DD",X"43",X"5F",X"96",X"47",X"90",X"43",X"BD",X"82",X"7B",X"10",X"83",X"02",X"80",X"2F",X"03",
		X"CC",X"02",X"80",X"10",X"83",X"FD",X"80",X"2E",X"03",X"CC",X"FD",X"80",X"DD",X"3F",X"5F",X"96",
		X"48",X"93",X"44",X"BD",X"82",X"7B",X"10",X"83",X"04",X"00",X"2F",X"03",X"CC",X"04",X"00",X"10",
		X"83",X"FC",X"00",X"2E",X"03",X"CC",X"FC",X"00",X"DD",X"41",X"DC",X"45",X"20",X"26",X"81",X"07",
		X"24",X"05",X"86",X"07",X"6C",X"C8",X"10",X"81",X"86",X"25",X"05",X"86",X"86",X"6C",X"C8",X"10",
		X"39",X"C1",X"39",X"24",X"05",X"C6",X"39",X"6C",X"C8",X"10",X"C1",X"D2",X"25",X"05",X"C6",X"D2",
		X"6C",X"C8",X"10",X"39",X"34",X"24",X"8D",X"38",X"E7",X"03",X"5F",X"96",X"43",X"ED",X"11",X"ED",
		X"15",X"96",X"44",X"A7",X"13",X"ED",X"17",X"DC",X"3F",X"ED",X"1C",X"DC",X"41",X"ED",X"1E",X"BD",
		X"D8",X"C6",X"31",X"84",X"BD",X"D6",X"8B",X"5D",X"B0",X"22",X"10",X"AF",X"07",X"AF",X"2A",X"10",
		X"9F",X"2A",X"35",X"A4",X"BD",X"5F",X"31",X"C6",X"05",X"BD",X"5D",X"BF",X"3D",X"48",X"20",X"03",
		X"BD",X"D7",X"50",X"A7",X"19",X"48",X"10",X"8E",X"00",X"00",X"10",X"AE",X"A6",X"10",X"AF",X"08",
		X"86",X"04",X"A7",X"03",X"39",X"96",X"BD",X"5F",X"A3",X"15",X"24",X"04",X"43",X"50",X"82",X"FF",
		X"58",X"49",X"DD",X"BF",X"96",X"BE",X"5F",X"A3",X"17",X"24",X"04",X"43",X"50",X"82",X"FF",X"D3",
		X"BF",X"24",X"03",X"CC",X"FF",X"FF",X"39",X"00",X"00",X"01",X"02",X"02",X"01",X"A6",X"4A",X"4C",
		X"81",X"06",X"26",X"01",X"4F",X"10",X"8E",X"89",X"57",X"E6",X"A6",X"E7",X"05",X"A7",X"4A",X"39",
		X"07",X"BB",X"07",X"50",X"83",X"50",X"83",X"BB",X"44",X"35",X"1A",X"50",X"20",X"26",X"1A",X"50",
		X"EC",X"47",X"FD",X"CA",X"04",X"EC",X"4B",X"4C",X"FD",X"CA",X"06",X"7F",X"CA",X"02",X"7F",X"CA",
		X"03",X"7F",X"CA",X"01",X"86",X"12",X"B7",X"CA",X"00",X"6A",X"4C",X"26",X"05",X"1C",X"AF",X"7E",
		X"D6",X"C5",X"6C",X"48",X"EC",X"47",X"FD",X"CA",X"04",X"EC",X"4B",X"FD",X"CA",X"06",X"EC",X"49",
		X"FD",X"CA",X"02",X"C6",X"0A",X"A6",X"4D",X"27",X"05",X"B7",X"CA",X"01",X"C6",X"1A",X"F7",X"CA",
		X"00",X"1C",X"AF",X"A6",X"4E",X"8E",X"89",X"7E",X"7E",X"D6",X"BC",X"00",X"01",X"02",X"01",X"BE",
		X"99",X"86",X"03",X"82",X"2A",X"03",X"BE",X"99",X"CE",X"AF",X"4B",X"EC",X"47",X"81",X"07",X"24",
		X"02",X"86",X"07",X"81",X"83",X"25",X"02",X"86",X"83",X"C1",X"39",X"24",X"02",X"C6",X"39",X"C1",
		X"D9",X"25",X"02",X"C6",X"D9",X"ED",X"47",X"86",X"19",X"A7",X"4A",X"1A",X"50",X"FC",X"2B",X"0D",
		X"FD",X"CA",X"06",X"EC",X"47",X"FD",X"CA",X"04",X"CC",X"2B",X"0F",X"FD",X"CA",X"02",X"A6",X"4A",
		X"44",X"C6",X"0A",X"24",X"07",X"86",X"11",X"B7",X"CA",X"01",X"C6",X"1A",X"F7",X"CA",X"00",X"1C",
		X"AF",X"6A",X"4A",X"27",X"08",X"86",X"05",X"8E",X"89",X"FB",X"7E",X"D6",X"BC",X"BD",X"5F",X"31",
		X"5F",X"A6",X"47",X"ED",X"11",X"ED",X"15",X"A6",X"48",X"A7",X"13",X"ED",X"17",X"AF",X"47",X"CC",
		X"2A",X"F9",X"ED",X"08",X"BD",X"D8",X"C6",X"86",X"80",X"A7",X"19",X"6F",X"0C",X"9F",X"2E",X"86",
		X"50",X"A7",X"49",X"6F",X"4A",X"AE",X"47",X"6A",X"49",X"27",X"57",X"10",X"AE",X"4B",X"A6",X"31",
		X"26",X"12",X"FC",X"99",X"86",X"10",X"BC",X"99",X"CE",X"27",X"03",X"FC",X"99",X"CE",X"ED",X"4B",
		X"A6",X"31",X"27",X"20",X"E6",X"15",X"A0",X"11",X"25",X"02",X"CB",X"06",X"C0",X"03",X"E7",X"15",
		X"E6",X"17",X"A6",X"33",X"8B",X"08",X"A0",X"13",X"25",X"02",X"CB",X"0C",X"C0",X"06",X"C1",X"DA",
		X"24",X"02",X"E7",X"17",X"6F",X"02",X"BD",X"8A",X"F1",X"26",X"06",X"8E",X"E6",X"67",X"BD",X"E6",
		X"AA",X"86",X"02",X"BD",X"D6",X"BA",X"AE",X"47",X"6C",X"02",X"86",X"04",X"8E",X"8A",X"55",X"7E",
		X"D6",X"BC",X"CC",X"8A",X"F1",X"ED",X"4B",X"CC",X"8A",X"D4",X"ED",X"4D",X"CC",X"85",X"1B",X"ED",
		X"C8",X"15",X"86",X"04",X"A7",X"C8",X"11",X"A6",X"11",X"81",X"45",X"86",X"03",X"24",X"01",X"40",
		X"5F",X"7E",X"85",X"DF",X"BD",X"D7",X"7D",X"0A",X"81",X"7E",X"D6",X"C5",X"A6",X"4A",X"4C",X"81",
		X"04",X"26",X"01",X"4F",X"AE",X"47",X"10",X"8E",X"89",X"CB",X"E6",X"A6",X"E7",X"05",X"A7",X"4A",
		X"39",X"10",X"AE",X"47",X"BE",X"99",X"86",X"8D",X"14",X"24",X"07",X"AF",X"4B",X"6F",X"22",X"7E",
		X"8B",X"21",X"BE",X"99",X"CE",X"8D",X"06",X"25",X"F2",X"AE",X"47",X"20",X"CF",X"A6",X"11",X"27",
		X"0E",X"A6",X"31",X"E6",X"33",X"C0",X"08",X"DD",X"BD",X"BD",X"89",X"35",X"81",X"0B",X"39",X"4F",
		X"39",X"A6",X"11",X"81",X"49",X"CC",X"8B",X"B6",X"24",X"03",X"CC",X"8B",X"87",X"10",X"8E",X"99",
		X"D9",X"BC",X"99",X"86",X"26",X"04",X"10",X"8E",X"99",X"91",X"ED",X"27",X"CC",X"02",X"00",X"ED",
		X"23",X"86",X"04",X"ED",X"25",X"10",X"AF",X"4B",X"AE",X"47",X"86",X"03",X"A7",X"05",X"8E",X"E6",
		X"75",X"BD",X"E6",X"AA",X"AE",X"4B",X"EC",X"07",X"27",X"19",X"10",X"AE",X"47",X"AE",X"15",X"A6",
		X"11",X"27",X"10",X"E6",X"13",X"CB",X"08",X"A7",X"35",X"E7",X"37",X"86",X"01",X"8E",X"8B",X"54",
		X"7E",X"D6",X"BC",X"CC",X"01",X"00",X"ED",X"03",X"86",X"02",X"ED",X"05",X"AE",X"47",X"BD",X"D7",
		X"7D",X"BD",X"DC",X"73",X"7E",X"8A",X"D7",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"08",
		X"08",X"08",X"08",X"08",X"08",X"00",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",X"04",
		X"04",X"04",X"04",X"04",X"00",X"86",X"0A",X"BD",X"D6",X"BA",X"86",X"20",X"A7",X"4D",X"6F",X"4C",
		X"6F",X"49",X"EE",X"47",X"C6",X"44",X"11",X"83",X"99",X"D9",X"26",X"02",X"C6",X"22",X"9E",X"1C",
		X"E7",X"0A",X"BD",X"EA",X"F2",X"2B",X"DE",X"BD",X"6B",X"F3",X"25",X"09",X"8E",X"E6",X"8C",X"BD",
		X"E6",X"AA",X"BD",X"8D",X"07",X"DE",X"1C",X"A7",X"4B",X"BD",X"8C",X"E9",X"86",X"01",X"BD",X"D6",
		X"BA",X"86",X"01",X"BD",X"D6",X"BA",X"AE",X"47",X"96",X"39",X"10",X"9E",X"58",X"8C",X"99",X"D9",
		X"26",X"04",X"44",X"10",X"9E",X"5C",X"44",X"25",X"61",X"96",X"39",X"85",X"40",X"26",X"32",X"1F",
		X"20",X"85",X"C0",X"26",X"55",X"C5",X"03",X"26",X"51",X"84",X"0F",X"8E",X"8D",X"27",X"A6",X"86",
		X"2B",X"1F",X"A1",X"4B",X"27",X"1B",X"8E",X"98",X"A3",X"E6",X"86",X"C1",X"04",X"24",X"12",X"8D",
		X"66",X"BD",X"8C",X"F8",X"8E",X"98",X"A8",X"E7",X"86",X"E6",X"4B",X"A7",X"4B",X"8D",X"7A",X"8D",
		X"67",X"6A",X"4C",X"2E",X"09",X"86",X"48",X"E6",X"4D",X"54",X"27",X"1E",X"ED",X"4C",X"6A",X"49",
		X"2E",X"16",X"A6",X"4D",X"A7",X"49",X"8E",X"98",X"A8",X"A6",X"4B",X"E6",X"86",X"6F",X"86",X"5D",
		X"26",X"04",X"E6",X"4A",X"E7",X"86",X"8D",X"40",X"20",X"87",X"8D",X"2B",X"A6",X"4B",X"BD",X"E9",
		X"72",X"C6",X"03",X"3D",X"8E",X"EA",X"F1",X"30",X"85",X"A6",X"15",X"E6",X"17",X"EE",X"47",X"BD",
		X"6B",X"F3",X"25",X"06",X"8E",X"E6",X"91",X"BD",X"E6",X"AA",X"BD",X"73",X"75",X"86",X"78",X"BD",
		X"D6",X"BA",X"8D",X"34",X"7E",X"D6",X"C5",X"34",X"06",X"A6",X"4B",X"8E",X"98",X"A8",X"E6",X"86",
		X"E7",X"61",X"6F",X"86",X"8D",X"04",X"35",X"86",X"A6",X"4B",X"8E",X"98",X"9E",X"E6",X"86",X"27",
		X"02",X"C6",X"02",X"8E",X"98",X"AD",X"E7",X"86",X"39",X"34",X"16",X"8E",X"98",X"A3",X"A6",X"4B",
		X"E6",X"86",X"CA",X"04",X"E7",X"86",X"35",X"96",X"34",X"16",X"8E",X"98",X"A3",X"A6",X"4B",X"E6",
		X"86",X"C4",X"FB",X"E7",X"86",X"35",X"96",X"D6",X"39",X"58",X"2B",X"1A",X"8E",X"D0",X"12",X"5F",
		X"30",X"03",X"EB",X"88",X"EE",X"8C",X"D0",X"2A",X"25",X"F6",X"C0",X"F2",X"27",X"08",X"D6",X"D2",
		X"26",X"04",X"0C",X"D2",X"0C",X"27",X"39",X"FF",X"01",X"03",X"FF",X"00",X"01",X"00",X"FF",X"02",
		X"02",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"2A",X"02",X"A7",X"03",X"39",X"2A",X"FD",X"BD",X"DC",
		X"73",X"A6",X"11",X"27",X"0A",X"E6",X"12",X"ED",X"15",X"A6",X"13",X"A7",X"17",X"6F",X"11",X"6C",
		X"02",X"39",X"8E",X"E6",X"99",X"BD",X"E6",X"AA",X"DE",X"1C",X"86",X"0A",X"A7",X"47",X"EE",X"4B",
		X"AE",X"55",X"A6",X"03",X"2A",X"03",X"7E",X"D6",X"C5",X"A6",X"02",X"26",X"F9",X"86",X"FF",X"A7",
		X"C8",X"23",X"6F",X"C8",X"24",X"BD",X"DF",X"C1",X"10",X"8E",X"8D",X"37",X"86",X"FF",X"8D",X"76",
		X"86",X"03",X"BD",X"D6",X"BA",X"EE",X"4B",X"BD",X"6B",X"F3",X"25",X"0E",X"96",X"39",X"2A",X"0F",
		X"48",X"2B",X"0C",X"C6",X"07",X"BD",X"37",X"B9",X"20",X"05",X"CC",X"74",X"AF",X"ED",X"4A",X"1A",
		X"F0",X"10",X"8E",X"8D",X"3C",X"8D",X"4F",X"AF",X"53",X"10",X"AE",X"55",X"A6",X"23",X"A7",X"03",
		X"4F",X"A7",X"C8",X"27",X"BD",X"8E",X"84",X"AE",X"55",X"86",X"02",X"BD",X"8E",X"84",X"AE",X"53",
		X"CC",X"1A",X"44",X"BD",X"8E",X"A4",X"AE",X"55",X"CC",X"0A",X"00",X"BD",X"8E",X"A4",X"1C",X"AF",
		X"86",X"03",X"BD",X"D6",X"BA",X"6A",X"47",X"27",X"3A",X"EE",X"4B",X"20",X"E1",X"AE",X"55",X"AD",
		X"A4",X"AE",X"59",X"AD",X"A4",X"AE",X"57",X"AD",X"A4",X"AE",X"5D",X"AD",X"A4",X"AE",X"5B",X"AD",
		X"A4",X"AE",X"53",X"AD",X"A4",X"39",X"AE",X"55",X"AD",X"A4",X"AE",X"59",X"AD",X"A4",X"AE",X"57",
		X"AD",X"A4",X"AE",X"5D",X"AD",X"A4",X"AE",X"5B",X"AD",X"A4",X"AE",X"53",X"2B",X"03",X"AE",X"C8",
		X"27",X"6E",X"A4",X"EE",X"4B",X"10",X"8E",X"36",X"AB",X"AE",X"55",X"BD",X"8F",X"06",X"AE",X"53",
		X"BD",X"8F",X"06",X"DE",X"1C",X"10",X"AF",X"49",X"86",X"07",X"BD",X"D6",X"BA",X"10",X"AE",X"49",
		X"EE",X"4B",X"A6",X"A4",X"26",X"E3",X"AE",X"55",X"CC",X"0E",X"10",X"8D",X"2D",X"AE",X"53",X"CC",
		X"07",X"0A",X"8D",X"26",X"BD",X"8E",X"C7",X"86",X"01",X"11",X"83",X"99",X"D9",X"26",X"01",X"4C",
		X"10",X"8E",X"8D",X"37",X"BD",X"8D",X"F6",X"1F",X"30",X"DE",X"1C",X"ED",X"47",X"96",X"39",X"43",
		X"84",X"03",X"27",X"03",X"7E",X"8B",X"EA",X"7E",X"D6",X"C5",X"1A",X"F0",X"FD",X"CA",X"06",X"A6",
		X"15",X"E6",X"17",X"FD",X"CA",X"04",X"FD",X"CA",X"02",X"7F",X"CA",X"01",X"86",X"12",X"B7",X"CA",
		X"00",X"1C",X"AF",X"39",X"A7",X"05",X"A7",X"04",X"C6",X"05",X"3D",X"E3",X"08",X"1F",X"02",X"EC",
		X"15",X"E3",X"22",X"ED",X"15",X"A6",X"17",X"AB",X"24",X"A7",X"17",X"10",X"AE",X"A4",X"31",X"22",
		X"10",X"AF",X"1A",X"39",X"34",X"07",X"6C",X"02",X"1A",X"F0",X"A6",X"15",X"E6",X"17",X"FD",X"CA",
		X"04",X"10",X"AE",X"1A",X"EC",X"3E",X"FD",X"CA",X"06",X"10",X"BF",X"CA",X"02",X"EC",X"61",X"F7",
		X"CA",X"01",X"B7",X"CA",X"00",X"35",X"87",X"96",X"39",X"11",X"83",X"99",X"D9",X"27",X"18",X"F6",
		X"99",X"11",X"26",X"31",X"85",X"01",X"26",X"2D",X"8A",X"01",X"97",X"39",X"7A",X"99",X"11",X"C6",
		X"5E",X"10",X"8E",X"2A",X"C0",X"20",X"16",X"F6",X"99",X"1A",X"26",X"19",X"85",X"02",X"26",X"15",
		X"8A",X"02",X"97",X"39",X"7A",X"99",X"1A",X"C6",X"5F",X"10",X"8E",X"56",X"C0",X"43",X"85",X"03",
		X"27",X"03",X"BD",X"69",X"5C",X"39",X"2B",X"05",X"A6",X"A0",X"26",X"FC",X"39",X"A6",X"15",X"27",
		X"F7",X"E6",X"17",X"1F",X"01",X"34",X"10",X"A6",X"A0",X"27",X"2B",X"84",X"0F",X"C6",X"11",X"3D",
		X"A6",X"3F",X"84",X"F0",X"44",X"44",X"44",X"44",X"26",X"06",X"6C",X"61",X"AE",X"E4",X"20",X"E7",
		X"27",X"E5",X"81",X"01",X"26",X"02",X"C4",X"F0",X"8C",X"90",X"00",X"24",X"DA",X"E7",X"84",X"30",
		X"89",X"01",X"00",X"4A",X"20",X"EA",X"35",X"90",X"86",X"02",X"A7",X"C8",X"25",X"6F",X"C8",X"27",
		X"86",X"04",X"A7",X"C8",X"26",X"BD",X"89",X"14",X"31",X"47",X"A6",X"C8",X"27",X"48",X"AF",X"A6",
		X"6F",X"11",X"BD",X"82",X"84",X"86",X"44",X"A7",X"0C",X"9F",X"2E",X"6C",X"C8",X"27",X"6A",X"C8",
		X"26",X"26",X"E2",X"86",X"01",X"BD",X"D6",X"BA",X"6A",X"C8",X"25",X"26",X"D3",X"31",X"47",X"86",
		X"08",X"97",X"3C",X"EC",X"C8",X"28",X"AE",X"A1",X"E7",X"17",X"E7",X"13",X"A7",X"15",X"A7",X"11",
		X"0A",X"3C",X"26",X"F2",X"31",X"47",X"C6",X"08",X"AE",X"A1",X"27",X"12",X"A6",X"11",X"26",X"0E",
		X"BD",X"D7",X"7D",X"A7",X"3F",X"A7",X"3E",X"6A",X"C8",X"27",X"10",X"27",X"47",X"17",X"5A",X"26",
		X"E7",X"86",X"03",X"8E",X"8F",X"94",X"7E",X"D6",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
