-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_1M is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_1M is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_1M_0 : RAMB16_S2
	generic map (
		INIT_00 => x"426F75C120B3AE2D610CE6B8A62B8AA216AA59C40B340279780B080B080B38A1",
		INIT_01 => x"2846219104D041351B28A60466058160710208E088339852426188515DCD422D",
		INIT_02 => x"8E2C7337587505A2C69898139E28D919E489A6492124927881159879C75D7F52",
		INIT_03 => x"864701678841055B28A6A1982F0862088E20F1F41626941D784A208822388709",
		INIT_04 => x"8223887D5E5EC75787B5361D79C61A622C41E71CF509234E7413BD8522F75218",
		INIT_05 => x"A8E4DAB3B2C2444B39822D66D2C5A2CEBB2AECE841607D87D04ED581A05AE218",
		INIT_06 => x"CECB3A1C758526549B5E89EB516549B505E418AC10CAECD824D0CA0ECD024D0C",
		INIT_07 => x"75D7135E5E8433B5D41C6988A171C1965881607C41251261098000000746637E",
		INIT_08 => x"A7E464A46424E4A4642415115D57111B445755C442D09AD3515E668926786045",
		INIT_09 => x"35ACD6B35ACD6B35ACD6B3506A298E20B86A298EDE4684E0426389144117A4A4",
		INIT_0A => x"390E4E5B38A283B2390E4E58E4E5B38A67A8E4488A688A499AA4E24E0A9ACD6B",
		INIT_0B => x"691B579D57BD875E10586208919281964B382240992CE588E39839AC66B293B6",
		INIT_0C => x"9AC49082388A2145D75454416F660663660400DAAAA9CAA4B882218AA2186062",
		INIT_0D => x"28209E19EA6892A788684E05E24E79C9B2A2C20432814CA063281D4A140524A0",
		INIT_0E => x"495909EB9DB9A7E2649514169C5C75361D4E228B5071A71078A26282089A0099",
		INIT_0F => x"000000000000000106A252265059E907E2A377CA5318A6A354555C65CDB0F59B",
		INIT_10 => x"6068F058161B681AC510410518535A730DDDD48024948659C0A6948E79452A45",
		INIT_11 => x"5A5DC57250812477708D5A494949494949858989898989898989B5898954AF41",
		INIT_12 => x"1A63F89144041341775C5C7FEB99471B585DD7151FA24514F1B5DE8FE8F1B515",
		INIT_13 => x"108292829180A846245065E04B56ED4E09AF1A6F3A5686595E62D858F2E05259",
		INIT_14 => x"14571F5E4182D3A5E6973A5EE7DAA415E59E21E0813954A0A42064A02A138B25",
		INIT_15 => x"0E7AE666E5E565E55AD532596972DE450C965A721861C8030C30046464646465",
		INIT_16 => x"146104905193938822188105904154115DF598198D98168D7D5D7D49F9D9F90A",
		INIT_17 => x"2548E657322473247ED55413C810557A4F2041F93C8105391904144124104124",
		INIT_18 => x"B2627141C413710F6BD0FE8D933F6F533F35BDA39B5507A25489A4E22415A261",
		INIT_19 => x"05498E0500D04D05BD5D9D9D9D9D9D9D9D9D9D9D9D9D929CFFD2552714172EEA",
		INIT_1A => x"62D9FC820209059388D4C235308D4E235388D4E235388D4D951D9514B579F049",
		INIT_1B => x"96AD616A9A61AAD616B4642D1FC8202094B9A249748925D224974A925D212674",
		INIT_1C => x"04906189522611049071441241C544124186DB254899516156EB896AD625AB5A",
		INIT_1D => x"5BA688208B45124907A62520458EA8A8E43992B88AA88A8B4B169B3A2CA8B391",
		INIT_1E => x"0000000000000000000004E2860822841241455C4BA68A2AAAAA2A861241C5DC",
		INIT_1F => x"2BAF7DC700000000000000000000000000000000000007F50000000000000000",
		INIT_20 => x"00000000004E6098E209FF73D8B4F4A1898115D516544144926542C50B08F005",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"5949B9191C9050B8141D04088B1B89058308A298220B9D909F929C5420821862",
		INIT_23 => x"8647461A411922E6758B9AF1D0942245198D68B95EDE989E98D8D8D08109B969",
		INIT_24 => x"898928908A0F02E4A046A19142E7A55787B2BD8A482E098225F1B4DA66224E93",
		INIT_25 => x"D517D22567545F4A999D517D22667545F4A959D517D22767545F4A91988AA2C8",
		INIT_26 => x"38604D7BD6BA465271B89058308A2982E7D26DE5DA4D655D517D2467545F69D9",
		INIT_27 => x"9EC9071270889EF1250B9EC98D05C64D241719E41146F739124EF7191E42E2BD",
		INIT_28 => x"98D8D88A7193490415C53D6798798D8D88A7191790468D5208B3127208A29A2B",
		INIT_29 => x"496269A25556DCCDEFD7896B95A94994A259535CB089389060B8E65051DA494C",
		INIT_2A => x"495055555555B51512696568D5B89054997896B95A949955055472BFD85572C9",
		INIT_2B => x"8815D55555557D454CD095458D034B8922415D5555550767D072567D07E7D07A",
		INIT_2C => x"BDF828790BD06641549EBE7AA5CBDDDD0A6415555555D4506625514E234EAE24",
		INIT_2D => x"02555FE6286C9CB9EA9CF0286C9CB9DA9559999F8284909DF8284909DF828590",
		INIT_2E => x"BAA4341E0A84A8A4341E0641E5126A90D07809EC8D489279A207862792820282",
		INIT_2F => x"04228A6279E78B116152C927BA781053B00A4228A628204228A6249AA4341A84",
		INIT_30 => x"A76524E4A76424E4A76724E4A76624E4A4642515E4A46424E4A4155927881E82",
		INIT_31 => x"208AC5A922022A38ED598E3A54638A19C2191097708207129C22A18308A298E4",
		INIT_32 => x"55C77429CDB36860EB212B0889097B09061A5A5546E3990504ED8E43B6063B0A",
		INIT_33 => x"A25B9265492094EED25581541DD06736CDA183AC84EC22242721906D75755550",
		INIT_34 => x"9A28DAE6B85A1608858ABAABAABA6C69E90A764E9F92A7A46BF0B82BB9A55789",
		INIT_35 => x"FC822AA0CEE0957D7A7A0A6B88A59AA3296698B996CA8668A36B8856698B8591",
		INIT_36 => x"54E42E08E555B94A9C723515539A08229A0821AA383BFFFC8239A0A18620BA1B",
		INIT_37 => x"B28A382849279188EE1818EE09555DF38A082A081A0954A08156954855472525",
		INIT_38 => x"00000000000000000000000000000000000000000000000000000000557BE49C",
		INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"01C7FE77D72C7ED3BCDE3DEF0000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1M_1 : RAMB16_S2
	generic map (
		INIT_00 => x"C039EBCF33918833CB000310C8330CC35C44484CC83248232921092119291847",
		INIT_01 => x"3CCC38384280C30D2138C300C33DCF30FB0810420C000C3300300D75DF22C033",
		INIT_02 => x"D03CF07CF2FB3C0B9FF20D318C3245ACE00CE3080C200C20CF100CF7CF7AF9CC",
		INIT_03 => x"E0E30F312E030D3138C3D30C86284320C4303BECBF0C8C3AFCCC320C0310CC50",
		INIT_04 => x"C8310CC3C8CACCF2329B7CBEF79F3FC83FCFDF32CD8CE6C65D31BFCC039EB330",
		INIT_05 => x"6A20F3918642888400C03AC046238C46091804ACCF38E7CF34C6ACCF73CC8330",
		INIT_06 => x"4A291B3CCF2E0E4C3B338CE931E0C3937E24B628B84624F66CF846620FE68F84",
		INIT_07 => x"223F37C8CA2C919BECF9FF20F38F210E10D334F3CF0042F300C0000006C03FC8",
		INIT_08 => x"DF9C9C5C5E5E1C1E1C1C8E32083084618C820C2114630F71E1CC302C032023C8",
		INIT_09 => x"3E2CF8A3E24F883E2CF8A3C9E759DE768D2368D24A9CC18014340E3404231CDC",
		INIT_0A => x"1A84C6791843E1191A84C6784C679184368C666142524268DE30834A30E24F88",
		INIT_0B => x"D028F203D2A71EBF33CCC320E106610E611843610D646604210719E46791A119",
		INIT_0C => x"3A2E90CA20C835D72CF8330BF6E22E13E12CC0F11115464E20C8320D67288CA2",
		INIT_0D => x"E8328808C302C0320DCC18000F072A6793944A0F938364E0F93836CC008330C3",
		INIT_0E => x"DF070763C7C73D433C8E0CBF717CDB7CB3C8320FB3E7FF3210C8330C20FEA20F",
		INIT_0F => x"00000000000000023C71C213C3CED301D1B0CCC4D9AC4F953221E1C707CE1DF1",
		INIT_10 => x"F3EE02FCFBA118F78EFBCF010CEAC49A33333E261CF8E1CF0A1CFC21CF333903",
		INIT_11 => x"06A32EF1E8C036CCD8D4C60707070707077307070707070707075307073466CB",
		INIT_12 => x"C6A0194CC910C1202A6C14C00CCC112D480A9B863037100252D44E8A6652D400",
		INIT_13 => x"4853EB52C850F9C8383123E08EEC73A30AC62A462AF19EF8C4333C28011CE208",
		INIT_14 => x"08C5300D90634BE5359099093B46800609847C603E4BD294FA1432D43E720FAF",
		INIT_15 => x"E3195D5D1D7D7D3CD93992001AB146AE64800641041050030C3002110033221B",
		INIT_16 => x"F1083C421796A10C4320CF1003C420F2089E88B84F84BC8F8717170317170763",
		INIT_17 => x"1308C38201142C962656020A040215A8281420A0A0500260703C480F0003C000",
		INIT_18 => x"D0F0D0FBCCCC10C1A50C1E50A040D020400373730D562D71F084E0C32F4031F8",
		INIT_19 => x"03C8C61340F1C72FFC800000000000000000000000000828050D800D0FB98B42",
		INIT_1A => x"D23CFE46A30A2FF848FE103F848FE013F800FE033F808FE3B3BF7F708C1700C3",
		INIT_1B => x"4AC08CAC081CAC08CADFDF2345446A30A23FE32B0224AC0852B0204AC08CADEC",
		INIT_1C => x"C07010C7C213C3C070100F01C0410F01C0439C1F084E23CC883F8CAC0852B020",
		INIT_1D => x"2B2328C288C0300723FE3C2808C83D8C6E20E3D142F242D1188EF11B646D91A3",
		INIT_1E => x"0000000000000000000008C28C28C18C01CCA3B22B2328418008038CC1C4A3F2",
		INIT_1F => x"04128338000000000000000000000000000000000000011B0000000000000000",
		INIT_20 => x"000000000084310CA10AFFB00C00AC038FC410CE1E4CC43000E0C2430908000B",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"171707838878392DCDB30E8DC49D4F73608CE30DC313E1717C7C703430883043",
		INIT_23 => x"9096D250CC5863BC40AEF30B307A334307CB19EF00327E7174BCB4BD00271717",
		INIT_24 => x"FF97C058F2EE2BBF002438300BBE1DE00092D7C70A4B82C430270F79C43FD034",
		INIT_25 => x"1D8C71BD1C7431C5F071D0C71BD1C7631C5F071D8C71BD1C7431C5F0718CA308",
		INIT_26 => x"5100174874A1F1D1D9F4F73608CE30C4F877C73C73C73E31D0C7BD1C7631DF07",
		INIT_27 => x"F3135E75F8C4F3275E0EF3134B6BCCC07C0F333C0014CC8C07D0CC8C03E4BF3C",
		INIT_28 => x"74BCBC23F3301F01971E4B7C76074B4BC23F3300F0104B9010CA75D88CE30D3E",
		INIT_29 => x"09A3084375DADCCDEFE41F40F40F40FBC3C7B63C560D9FFDC0D56975E5B7D721",
		INIT_2A => x"D7B40D75830D4B1133CF1D04B6BCF4352F42F41F41F41F3682ADB1C02E2AB1C7",
		INIT_2B => x"C50C0DDD603362C04298EEC44B626BCFB1D0C0DDD6030D3C30D3EEFC0D3C30D3",
		INIT_2C => x"EBA237FFEEB633C034FC43D13EC53333A33C075603372C00D03BB12892E9AF3E",
		INIT_2D => x"E380389637F0FE4F74FA2637F0FE4F44F7350CF2237CFCEBA237CFEEB2237CFC",
		INIT_2E => x"0F433CBF47A90D423CBF470BF6A43904F2FD1CACCF30E482033EEA72A32363A3",
		INIT_2F => x"98338C3100000D91C4E44E68198870206E8E8338C33CB98338C3191C403CBF29",
		INIT_30 => x"1E1C1C9C9E9C9C1C1E1F1C9C9E9F9E1E1F1D1D8D5D5C5C5C1C1C8E82020CFBCF",
		INIT_31 => x"0BCAE42D03C3280CA5E76F3978DBCE176739717AD9CE5C7076F287608CE30C1C",
		INIT_32 => x"BBC2EDBE07C1FA14FC0A3A0E8707809E00853137A6B2A3230C4446A1118B1B0D",
		INIT_33 => x"0F42D0F862CB6431DA63EEEC0BB6F81F07E853F028E83A1C1E09E000531378FB",
		INIT_34 => x"CE190CF18A388C19A3868F9B1E8B547A251E8543A050E8943800D468BCE5A41D",
		INIT_35 => x"BB4611CB2311A033202A8E33D6F38C34ACE30D89CEA323386433DE8E30D8A3B8",
		INIT_36 => x"5AFE388CE6340F40FFF92E0DE00C84600C84600C858FBBB84600C0D8C4313F0F",
		INIT_37 => x"500C9F08CCC3800FA3030BAF19560C918C8D0E8D0C8FFC59C00CFBDE3ADB1C27",
		INIT_38 => x"000000000000000000000000000000000000000000000000000000008034DB0C",
		INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"090871071C61830090A1CB240000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1M_2 : RAMB16_S2
	generic map (
		INIT_00 => x"0F32048CB031C3330800333CC330CC331088CC08482B0B1F1C230C233C233C08",
		INIT_01 => x"32033182AF0D20B0132CB3303332CC3B1C033CF2CC00CC810F30CC4100120F33",
		INIT_02 => x"C7360810C21880B73000CC02CB31809CB2ECD32CBCB3CB2CC000A228A1C1220B",
		INIT_03 => x"C6094C333F3480132CB3C0CCB42C730CCF331C72431124C1220330CC333CCC1C",
		INIT_04 => x"C333CCC307C760C1F1C01086283080033620A281A08CB20B0002D820F320430C",
		INIT_05 => x"B9040332C4CF00000CCF3307CF10C0CB132C4C320C300821800B10CCB30C330C",
		INIT_06 => x"C3031C8A0C20106440915CB091024429200C410C42CB08010802CB500050002C",
		INIT_07 => x"18318107C720B1C06203000CC80013C32CC030200030EA083CC0000000033100",
		INIT_08 => x"37343434373734353434A4E106044D03384142138CC0CC82090B32DCB31CF004",
		INIT_09 => x"000800200080020004001034C330C8320C8310C4C706E8628731CCE0402B7434",
		INIT_0A => x"1C43C3330CB351E41E43C3303C3130CB304C7520B330B320CC3C33C30CC0C003",
		INIT_0B => x"0A3CC2F332C82048830C330CC3CF13C3032F331CCCCCB30872CB2C3CF032C1E4",
		INIT_0C => x"8E1388CB3CCF310420C082243103102001100002222011390CCF33CC533CFCF2",
		INIT_0D => x"E232C73CB32DCB32CC6E8628FF672CD032C0CF41B2F0ACB82B2D010A084810E3",
		INIT_0E => x"4D0D0D03CDC9244334E4A24300460010830F33CD880C02812CC3338E2CCE12CC",
		INIT_0F => x"000000000000000032330B01E32C362732A6660A48FCA4049283434D8DE134D3",
		INIT_10 => x"332C090CCB331CCB20C30020220007C44999912314F6314FA714FAB14F1B0009",
		INIT_11 => x"8704DD4348C9BDE648D2472D0D2D0D2D0D590D2D0D2D0D2D0D2D492D0D98A124",
		INIT_12 => x"C7367405D404E0E4A28F0E169C01084CF928A3C3867024A2C4CFCBD6D2C4CCD3",
		INIT_13 => x"C4CAC6C9D4C8F3073083009BC884C0A32C481C081C0330000732210DA30ED04A",
		INIT_14 => x"545686634123CBD90024B1799507081C52473C72FC003172B13235B23CC1CF40",
		INIT_15 => x"231C3434373737366134B04E1C5107DD2C1387FF3CF3FC030C30077777666661",
		INIT_16 => x"030E0002A1A182CF333CC0106004380106200C40800440000DCDCDC40D0D0D23",
		INIT_17 => x"032C330B6380884088E0CBBC8C82A30CF2301223C8C0481A1A00408010200418",
		INIT_18 => x"C371024438C281DBD1ADB112F6FB06B6FB481490CD9090B332C0783323E2F31E",
		INIT_19 => x"4900C759100A2890FC88888888888888888888888888880DAC240610244CFB0E",
		INIT_1A => x"020E0187233C90C81002040081C02070081C020600818020440CC88881888304",
		INIT_1B => x"0B10BCB10B2CB10BCB03212060287233C2DCDB2CC2C0B30B02CC2C0B30BCB211",
		INIT_1C => x"14C112CCCB01EE04C112F893044BF853044BBE332C0782040B716CB10B02C42C",
		INIT_1D => x"2C030C618581E14C01C5BCB580C3334C710CC330B330B33F3C43132C8CB331CE",
		INIT_1E => x"000000000000000000000020820820B8130058812CC30CE28E28E1B8530478C1",
		INIT_1F => x"0820430800000000000000000000000000000000000003000000000000000000",
		INIT_20 => x"00000000000F33CD82CC00250D4DA5444DC0286410678018910A5CDC733C0010",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"0F0F0F0820F0B1CCA779348DC28C8D29D08CB2CCB31FCCDCD8D8D09633C30C73",
		INIT_23 => x"8E4D8E398139D735464CD537B0F2330B0D0154CD7100D8D0D0101413820F0F0F",
		INIT_24 => x"CDCD3D48CF207334E0833082633436C3C3C4C3332C730CC7370D40D055734E63",
		INIT_25 => x"60ACD4343581B354D0D60ECD8343580B364D0D60ECDC343580B374D0D77D5B45",
		INIT_26 => x"38E08D0CD0E3634378C8D29D08CB2CC7F0F34F34F34F34B60ACD343581B34D0D",
		INIT_27 => x"D71060D50BF8D70D50DCD710C13F718D2421C624234E70FC234E70FC2347338E",
		INIT_28 => x"DC181323DC63490B4D35362495CDC181323DC6349098C1031CE4D5348CB2CDFC",
		INIT_29 => x"2D832CB3B260840048C0CD0CD0CD0CD0E2CB75B443CCCCD368C8F0D35362495C",
		INIT_2A => x"C3506696292D0101C101058C163CD092CF2CF2CF2CF2CFB840A0A2EA8702808B",
		INIT_2B => x"002CA6E5019B71414308F1C1C32063CF0042CA6E5099373E9373D5B5373E9373",
		INIT_2C => x"C142373F2C1A3341B84063C13D44BBBB33372B9019B71413503C7070B0F18F3C",
		INIT_2D => x"3B06BD1C3738400F00F5423738400F00FBB70CD02372F2C102372F2C142370F2",
		INIT_2E => x"CD4D02436790CD4D024367E43C433134090D9CB3002CC30C3332D172C3333B33",
		INIT_2F => x"CE32CB305DF7CC5132438430E10C8428B68FE32CB31AFCE32CB300CF4E024350",
		INIT_30 => x"BEBFBC7E7E7F7E7C7E7E7E3E3E3E3F3F3C3D3C6D353434343434A40C32CCCBAF",
		INIT_31 => x"C8CB90CC33272C8CB3502F2CD70BCB0DB32CD0D50CCB34D0D3F2CDD08CB2CCBC",
		INIT_32 => x"75E6E4CF8FE37102FDCB2D8F0F0D449F01A7B7991132DC2930380311E0371D8E",
		INIT_33 => x"330FC3B01F07B2320709D1D49B933E3F8DC40BF72CB63C3C37C9F0127B799274",
		INIT_34 => x"CB150BF1672F4B5572C5C4050DC00236008D80235008D4023608C8763CB400DC",
		INIT_35 => x"30B31CC7232CCC4C1C1C8F2FD372CB35CCB2CD64CB63632C542FDFCB2CD672C8",
		INIT_36 => x"82F23D8C3C91CD1CDA08042643CC8B33CC8B33CC408F3333B30CC8C4C330FC8F",
		INIT_37 => x"41CCCF1F803421CD131F1D0F1E4CC4DFD0408C508D8FFD0CC0A4D107920A2CB9",
		INIT_38 => x"00000000000000000000000000000000000000000000000000000000318EF4E4",
		INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"051041C6186187104041C6180000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_1M_3 : RAMB16_S2
	generic map (
		INIT_00 => x"E405DF8F86E82404DF3E0090240902405DDD59994F4113A0A04EA04E904E901F",
		INIT_01 => x"04E80904C930C34F7E924032803C0F04DF28924800F800F0240A0176DF05E407",
		INIT_02 => x"2407DB4D37DF4E807DF9017828000C2E8A0137A2828A28A00F0284CF3DF7E5E8",
		INIT_03 => x"24130F07DDC30F7E92404A020B8280A02407DF7D303F4CF7E4E80A0280901390",
		INIT_04 => x"28090134E8287D3A0A1F4DF7CF7D37E407D33CF03C0E84E06D781F4E805DF0A0",
		INIT_05 => x"0038F7E813A4CCCF802404D3A80B1FA07E81FA84CF04D74DF5E07C0F03C240A0",
		INIT_06 => x"A87E8133D37F3FCCFF35CE8F33FCCFE36F34F034F0A034F034F0A0038F038F0A",
		INIT_07 => x"A34DF4E8287C281F7D37DF9013DF092CB01705E7CF0284D39000000004E807DB",
		INIT_08 => x"0F0E0C0C0D0D0C0C0C0E0FB028B0285EEC0A2C0A13BA0133F4E80A0280A243C0",
		INIT_09 => x"3F3CFCF3F3CFCF3F3CFCF3C1F37CDF37CDF37CDFA8E4F243240903B800830C0C",
		INIT_0A => x"8028285EA200080B8028285E8285EA2004CE0C5CE04CE05CD33E80E8A033CFCF",
		INIT_0B => x"D0913A37FA177DF933C280A03928092C7E82000801BA06DE080C81FA47E8380B",
		INIT_0C => x"3C0F00EC902405DB5DFCF01306CF3CF3CE3C30F7777755489024090133924243",
		INIT_0D => x"C03B289280A0280A024F24328003A3C6E91FA44F2903CA40F29035E4000F0249",
		INIT_0E => x"C703036FC7471DB31E4F4D306D77DF4DF4E40901F4DF7CF0A0240924B03C0B03",
		INIT_0F => x"00000000000000033CD3E80303C307020B30CC6CC026CD0A3830F1C707401C71",
		INIT_10 => x"03C1B4C0F05EA0F84D77CF1204F5E843033330002C7002C7002C7002C7A30083",
		INIT_11 => x"28DBC0C0C0C00C0CC0E0E8030333332323832313130303333323A33303FEC6D3",
		INIT_12 => x"28F01028C002C1F3F3CF3C000428A181FCFCF3CF00108204981F68C040981E08",
		INIT_13 => x"0000C001C100D6E00CF217B265DF9B4381F7813781F46DF5E809703C000C0020",
		INIT_14 => x"300F00F0000343CF0060263D11A8600DF6E8328801F7C0403000700035B8021F",
		INIT_15 => x"03A00C0C0F1F1F1FF7C02020A310A8C0080828FF3CF3FC030C3009999999999F",
		INIT_16 => x"F3243C483939380200900F02C3C0A0F0285F3CF3CF38F34FC7C7C7CF03030303",
		INIT_17 => x"00A280FF00481F481FBFFF2400083FDB9000206E40008393933C080F02C3C0B0",
		INIT_18 => x"2803E8DB6C0628C1428C142470110A3011901F4A01FF4CD3CA00C2803D4A13F0",
		INIT_19 => x"D34CE0C330F4D34C3C44444444444444444444444444443C0680FF3E8DB684A1",
		INIT_1A => x"63D400E003934C173CF5CF3D738F5CE3D738F5CE3D738F5D55511110F40D73CF",
		INIT_1B => x"E84E8284E83284E82847773DC01E00393A01B3A1BA0E86E83A1BA0E86E828666",
		INIT_1C => x"90F0384F28030BA0F038EE83C0C3EE83C0C1343CA00C33C0E804CE84E83A13A0",
		INIT_1D => x"A13392CB2DC0BB0F001F328F0C2806CE00A0306CE06CE06EA02C6E81BA06E83B",
		INIT_1E => x"000000000000000000000ECB2CB2CB2EC3C0F170A13392492492492E43C0E1B0",
		INIT_1F => x"1F7DF4D300000000000000000000000000000000000005DF0000000000000000",
		INIT_20 => x"0000000000E40901778300E5C17C0D75CB40B28F3F4EC0A2C3F0D3934E90F013",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"03030380403838224F031C0C010CC793C00E490240A33434303839303928A280",
		INIT_23 => x"2425E491C091F31D37DC74F03030348303CF7EC74D703C303CF8FCFA00030303",
		INIT_24 => x"C743A0C0E807071E83200800071C0FFA2A181803A208822804C35C72D371E479",
		INIT_25 => x"4E0C731D0D3831CC7434E0C731D0D3831CC7434E0C731D0D3831CC7436CDF34C",
		INIT_26 => x"924007807800E0C0D0CC793C00E49028CC71C71C71C71FF4E0C71D0D3831C743",
		INIT_27 => x"74DF4C36C0CC74C36C0C74DFCF093DC41C04F71C01243C1C81E43C1C81E08A0C",
		INIT_28 => x"38FCF0034F710700071C971C7C43CFCF0034F71070174FE0A03036F00E49003C",
		INIT_29 => x"A173A280FFFC840048F807807807807E81C7373429000C70C0CE4C71C971C704",
		INIT_2A => x"C7303FFFFFFD730173C71D74F5FC7A3A07A07A07A07A07FCE00510400C001040",
		INIT_2B => x"028E8FFFFFFF6CC07CC0D0C0CF077FC701E8E8FFFFFF1D1C31D1CDFC1D1C31D1",
		INIT_2C => x"4FF037F704F031C0FCF641D91C423333031D0FFFFFF7CC01D334303C13CD3F1C",
		INIT_2D => x"07FFF7DF37D0F4C74C70F037D0F4C74C7FF7CC7F037F704FF037C704FF037C70",
		INIT_2E => x"00073D30030A00073D3003D30D28001CF4C00E810FA028A2803C133A300F0B0B",
		INIT_2F => x"4C392400A28B0303D4E80E8A03A0F030D00DC392400C74C392400A00073D300A",
		INIT_30 => x"0C0E0E0D0C0E0D0E0C0E0D0D0C0E0D0D0C0C0E0C0C0C0C0C0C0E0F820A00F8C3",
		INIT_31 => x"00E009024003810E00DB0F8034C3E00343803037C0E00C30303803C00E49020E",
		INIT_32 => x"33F0CC0D0741D000F402800D03036C0D034A3A3FDB381F833E80E808030B800C",
		INIT_33 => x"4890248F8103D03360FF80CC0330341D074003D00A00340C0C00D0388383FFE0",
		INIT_34 => x"E807E8C07EA32887EA017006CD700035C00D70035C00D70037C0CE07FE8FF932",
		INIT_35 => x"CCE0800003383FDFA2A00DA3003A28000E8A007CE80303A01FA300A8A007EA00",
		INIT_36 => x"F4F4350E8FF8078073C13E0FF9002E09001E09000C0CCCCCE0A000C0280A300C",
		INIT_37 => x"2A000CA2C0A00A0133A0A13FA3FFF65A50100C000C0C0000C0FC735C3051028F",
		INIT_38 => x"00000000000000000000000000000000000000000000000000000000FFC0C284",
		INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"04D34D37DB7DF4D34C7DF5DF0000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
