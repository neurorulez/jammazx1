-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "281E03C01F802D5E3D542D5E07BC003C00782D5E281F3F550BC017D41C2D0B58";
    attribute INIT_01 of inst : label is "3C003C003C003D553C2D3D781E0A0B5E3C0F3D5E1E2D3C0F3C0F05783D0C255E";
    attribute INIT_02 of inst : label is "0000000000000000FFFF2FF8FFFF2FF807D0000007D000000140000001400000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0618000006180000000006000000000001FF0000FF000000000500AF4000FF40";
    attribute INIT_05 of inst : label is "00000000F000E0000F000BFFF000BFFFF0F0F0F0F0F0F0F005550FFFF00FF00F";
    attribute INIT_06 of inst : label is "007802803F540AA82AAD0AA81E3C002801F40AA8017E2AAA03C02AA83C0F02A0";
    attribute INIT_07 of inst : label is "C000D555C000C000000355570003000301500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C0002A83D5428003D542AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA803C02AA83D5F280A";
    attribute INIT_0A of inst : label is "3DDF08083D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "80000000E86A80AAEA4A8000C683255803E0080001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "002A0000003F003FAAAA0000F400FFFF2AAA00003FC03FFF0002000000000001";
    attribute INIT_0D of inst : label is "00000000000000002AAA00000000000702AA000003FD03FFAAAA00000000FFFF";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0008000A30C3A828330C80A0030C0802AA4C2A02090C2A02030C0A8200000000";
    attribute INIT_11 of inst : label is "000000003000800030CC0A02A4C3A028000A000290C3A0280000000218C3A828";
    attribute INIT_12 of inst : label is "002D000A5E00A8000FFC003001001300000200000C006000002F000AD6003000";
    attribute INIT_13 of inst : label is "0FF000A0F000000000153FF40000FC002FEF6800F80000000000002F3DFCFBE0";
    attribute INIT_14 of inst : label is "002900026800800001410296C140968000000000080000000001000080000000";
    attribute INIT_15 of inst : label is "35AA0000AA5C0000000110005400000400B300003800000000000F5C0000D7C0";
    attribute INIT_16 of inst : label is "000000000000000000000000000000007F5CFFFC3FFD3FFF0000FFD0000007FF";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "C240C00001830003C2400A55018355A0C300C30000C300C33015C300540C00C3";
    attribute INIT_1B of inst : label is "000000000000000000005555000055555555000055550000C015C300540300C3";
    attribute INIT_1C of inst : label is "000000C0000003005555000055550000000030000000000C0A55000055A00000";
    attribute INIT_1D of inst : label is "00D5000057000000000000C100004300002500005800000000C000C003000300";
    attribute INIT_1E of inst : label is "000000C0000003000180000002400000540000C000150300000055570000D555";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000540000C0001503000025000058000000";
    attribute INIT_20 of inst : label is "002D00300FFC000A5E0013000100A8000008002800BF00013000C00058008000";
    attribute INIT_21 of inst : label is "0FF02FF4001500A0F000FC00000000002FEF002F00006A00F800FBE03DFC0000";
    attribute INIT_22 of inst : label is "002902960141000268009680C140800000000000000100000800000080000000";
    attribute INIT_23 of inst : label is "35AA100000010000AA5C00045400000000B30F5C000000003800D7C000000000";
    attribute INIT_24 of inst : label is "3FFF10FC01FF0A02FFFC3FF4FF4080A03FFF10FC01FF2028FFFC3FF4FF402808";
    attribute INIT_25 of inst : label is "00FF000700000A80FF00D740000002A00FFF000700002A00F800D74000002A00";
    attribute INIT_26 of inst : label is "000000000000AAAA000000000000AAA0000000000000AAAA054000000000AAA0";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000FE00FFFC000000000000000000003FFF07FF0007FFFFFFFEFFFFFFFFFE00";
    attribute INIT_29 of inst : label is "FFF4F4000000A8000000000000000000002F0FFFBFFF0000FFFFFFFFFFF400AA";
    attribute INIT_2A of inst : label is "FFFEFFFFFFFF80008000FF40400000003FFF07FF0007FFFFFFFFFFFFFFFFFFFE";
    attribute INIT_2B of inst : label is "FFFFFFFFFFD4A800E000FFC000000000002F0FFFBFFF0000FFFFFFFFFFFF00AA";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFF0FF404000FFFC3FFF07FF0007FFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFA800E000FFC0FFF80000002F0FFFBFFF0000FFFFFFFFFFFF00AA";
    attribute INIT_2E of inst : label is "396907FF00000A006960FF40BD000280396907FF000000806960FF40BF800800";
    attribute INIT_2F of inst : label is "58D50C8300000000262633330000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "3FFF1FFC01FF0A02FFFC3F04FF4080A03FFF1FFC01FF2028FFFC3F04FF402808";
    attribute INIT_31 of inst : label is "3FFF1FFF01FF0A02FFFCFFF4FF4080A03FFF1FFF01FF2028FFFCFFF4FF402808";
    attribute INIT_32 of inst : label is "3FFF10FC01FF0A02FFFC3FF4FF4080A03FFF10FC01FF2028FFFC3FF4FF402808";
    attribute INIT_33 of inst : label is "3FFF1FFF01AF0A02FFFCFFF4FA4080A03FFF1FFF01AF2028FFFCFFF4FA402808";
    attribute INIT_34 of inst : label is "00C206C30000000058960CC3000000001D5220330000000058960CC300000000";
    attribute INIT_35 of inst : label is "C962CC230000000058960CC300000000256230330000000058960CC300000000";
    attribute INIT_36 of inst : label is "00003FE007FF000000002FF0FF4000000FFF3FE007FF000040000000E0000000";
    attribute INIT_37 of inst : label is "0FE03FFE07FF00002FC0FFF0FF4000000FFF3FFE07FF0000FFC08000FF400000";
    attribute INIT_38 of inst : label is "000000000000000000000000000000000FFF3FFF07FF0000FFC0FFF0FF400000";
    attribute INIT_39 of inst : label is "3FFF1FC701FF2028FD00FC74FF4020003FFF1FFF010F2028FD00FFF4F0402000";
    attribute INIT_3A of inst : label is "00A8BFFD10000000A800FFF80010000002BF3FF414000000FA007FF000500000";
    attribute INIT_3B of inst : label is "0AA0FF55000000002A8057FC0000000000A8FFF500000000A8007FFC00000000";
    attribute INIT_3C of inst : label is "BFFE000500000000FFF84000000000002BFE005500000000FFA0540000000000";
    attribute INIT_3D of inst : label is "007F000100000000F40000000000000017FF000100000000FF50000000000000";
    attribute INIT_3E of inst : label is "00030001000000000000000000000000000F000100000000C000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000400240000000000900080000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407E8014003C001503C0F";
    attribute INIT_01 of inst : label is "15553EA815553EA815503C0F01543C0015543EAD01503D5F05540AAF05501AF5";
    attribute INIT_02 of inst : label is "00000000000000001FF4FFFF1FF4FFFF00000BE000000BE00000028000000280";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0F3C00000F3C000000000F0000000000000500AFFFC0E800000001FF0000FD00";
    attribute INIT_05 of inst : label is "00000000D000F00007FF0F007FFFF000FFD0F0F0D0FFF0F003FF0FAAFFFDF00F";
    attribute INIT_06 of inst : label is "3EAF03C007E83C0F3EA8140F01FC2ABE0ABE140F1EAD1F8007C003C006B42F0E";
    attribute INIT_07 of inst : label is "C000C000EAAAC00000030003AAAB000300000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D2F3EAA3C003EAA3C003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F2BE803C03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "000040000000C02A0000EA001AA4C94300FC02002ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "003F00000000003FFFFF00000000FF503FFF000000003FF40003000000000000";
    attribute INIT_0D of inst : label is "000000000000000001FF00000000000003FF0000000003FFFFFF00000000D400";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "00060001706930C391A4330CEAC60C0CEA8640CCAB8640CC0706030C00000000";
    attribute INIT_11 of inst : label is "00000000900030001A4630CCA8690CC3000E0004B8690CC3000A0004A46980C3";
    attribute INIT_12 of inst : label is "003000006300C00001500BF000000300000600094C008C000005000154001800";
    attribute INIT_13 of inst : label is "0FF80BF0700020000000154B0000F4001E5F1F7AA78000000000001E05055F98";
    attribute INIT_14 of inst : label is "00C7000CC700700000050C7C58007C7000000000030000000000000200000000";
    attribute INIT_15 of inst : label is "2F550AFF55F8FFA00000000F0000F8000BFB0003BF80000000000C00000000C0";
    attribute INIT_16 of inst : label is "00000000000000003E2C000038BC0000BFA0FFFC0FFE3FFF0000F5000000005F";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "C300C02A00C3A803C300302A00C3A80CC300C30000C300C305AAC180AA500243";
    attribute INIT_1B of inst : label is "0000AAAA0000AAAA0000AAAA0000AAAAAAAA0000AAAA0000C000C18000030243";
    attribute INIT_1C of inst : label is "0000001A0000A4000000000000000000000005AA0000AA5030000000000C0000";
    attribute INIT_1D of inst : label is "00C2000083000000000000EA0000AB0000C000000300000000C000C003000300";
    attribute INIT_1E of inst : label is "0000001A0000A40000C0A8000300002A00000240000001800000AAAB0000EAAA";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000AAAA0240AAAA018000C0000003000000";
    attribute INIT_20 of inst : label is "00300BF001500000630003000000C00000190004001500269000600050003000";
    attribute INIT_21 of inst : label is "0FF8154B00000BF07000F400000020001E5F001E00001F7AA7805F9805050000";
    attribute INIT_22 of inst : label is "00C70C7C0005000CC7007C705800700000000002000000000300000000000000";
    attribute INIT_23 of inst : label is "2F55000F00000AFF55F8F8000000FFA00BFB0C0000000003BF8000C000000000";
    attribute INIT_24 of inst : label is "3FFF0FFF00053FEFFFFCFFF05000FBFC3FFF0FFF00053EFEFFFCFFF05000BFBC";
    attribute INIT_25 of inst : label is "001F000100000FFFFF00E3800000FFF001FF000100003FFFFE00E3800000FF00";
    attribute INIT_26 of inst : label is "0000000000001F550000000000005FF40000000000001FD7000000000000FFF4";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "E000FFE0FD50000000000000000000001FFF007F0000FFFFFFFFFFFF15FFFFE0";
    attribute INIT_29 of inst : label is "FF4040000000FFF8000000000000000002FF3FFFFFFF0002FFFFFFFFFF40BFFF";
    attribute INIT_2A of inst : label is "FFFFFFFFFD50FE80FE80F400000000001FFF007F0000FFFFFFFFFFFF15FFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFD400FFFAFE00D4000000000002FF3FFFFFFF0002FFFFFFFFFFFFBFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFD50FFFFFFD0F4000000FFFC1FFF007F0000FFFFFFFFFFFF15FFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFAFE00FFF0FFFC000002FF3FFFFFFF0002FFFFFFFFFFFFBFFF";
    attribute INIT_2E of inst : label is "1FDF001500002FFADFD052005000BFE01FDF001500002FEADFD050001400AFE0";
    attribute INIT_2F of inst : label is "A418501400000000333304040000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "3FFF0FFF00053FEFFFFCFFF05000FBFC3FFF0FFF00053EFEFFFCFFF05000BFBC";
    attribute INIT_31 of inst : label is "3F0F0FFF00053FEFF0FCFFF05000FBFC3F0F0FFF00053EFEF0FCFFF05000BFBC";
    attribute INIT_32 of inst : label is "3FFF0FFF00053FEFFFFCFFF05000FBFC3FFF0FFF00053EFEFFFCFFF05000BFBC";
    attribute INIT_33 of inst : label is "3FFF0F5F00053FEFFFFCF5F05000FBFC3FFF0F5F00053EFEFFFCF5F05000BFBC";
    attribute INIT_34 of inst : label is "75D30040000000000CC350140000000001830540000000000CC3501400000000";
    attribute INIT_35 of inst : label is "CE934140000000000CC35014000000001A930540000000000CC3501400000000";
    attribute INIT_36 of inst : label is "3E001FFE0015000002F0FFD0500000003FF41FFE001502BF000000005000F000";
    attribute INIT_37 of inst : label is "3FF81FFF00150280BFF0FFD050000A003FFF1FFF001502BFD400FE805000FA00";
    attribute INIT_38 of inst : label is "000000000000000000000000000000003FFF1FFF001502BFFFF0FFD05000FA00";
    attribute INIT_39 of inst : label is "3FFF0FFF00053EFEFF80FFF05000B8003FFF0FFF00053EFEFF80FFF05000B800";
    attribute INIT_3A of inst : label is "2FFFFF4000000000FFE007FC000000000FFF3F4000000000FFC007F000000000";
    attribute INIT_3B of inst : label is "BFFF000000000000FFF80000000000002FFF540000000000FFE0005400000000";
    attribute INIT_3C of inst : label is "15FF0000000002A0FD50000000002A00FFFF000000000000FFFC000000000000";
    attribute INIT_3D of inst : label is "001F0000000002FED00000000000FE00005F000000002FF8D40000000000BFE0";
    attribute INIT_3E of inst : label is "00030000000000030000000000000000000700000000002E400000000000E000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000005000024000002180280610000009000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "281E03C01F802D5E3D542D5E07BC003C00782D5E281F3F550BC017D41C2D0B58";
    attribute INIT_01 of inst : label is "3C003C003C003D553C2D3D781E0A0B5E3C0F3D5E1E2D3C0F3C0F05783D0C255E";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0618000006180000000006000000000001FF0000FF000000000500AF4000FF40";
    attribute INIT_05 of inst : label is "00000000F000E0000F000BFFF000BFFFF0F0F0F0F0F0F0F005550FFFF00FF00F";
    attribute INIT_06 of inst : label is "007802803F540AA82AAD0AA81E3C002801F40AA8017E2AAA03C02AA83C0F02A0";
    attribute INIT_07 of inst : label is "C000D555C000C000000355570003000301500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C0002A83D5428003D542AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA803C02AA83D5F280A";
    attribute INIT_0A of inst : label is "3DDF08083D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "80000000E86A80AAEA4A8000C683255803E0080001F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "002A0000003F003FAAAA0000F400FFFF2AAA00003FC03FFF0000000000000000";
    attribute INIT_0D of inst : label is "00000000000000002AA800000000000702AA000003FD03FFAAAA00000000FFFF";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0008000A30C3A828330C80A0030C0802AA4C2A02090C2A02030C0A8200000000";
    attribute INIT_11 of inst : label is "000000003000800030CC0A02A4C3A028000A000290C3A0280000000218C3A828";
    attribute INIT_12 of inst : label is "002F000AFE00A8000010003F0100FF00003D002FF3009E00001000350100CF00";
    attribute INIT_13 of inst : label is "0FFF00AAFFF00000001F3FFFFFD0FFF837FF6800F8000000000101F7F3FCFFE0";
    attribute INIT_14 of inst : label is "0000000000000000000000008000000003FF0000F7C0000001510FFF9500FFF0";
    attribute INIT_15 of inst : label is "3FFF0000FFFC000000003FFF0000FFFC0003000000000000000103FF0000FF00";
    attribute INIT_16 of inst : label is "00000000000000000000000000000000F4BCFFFC3FD23FFF0000FE90000007FA";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000AAAA0000AAAA000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "FF40FFFF01FFFFFFFF400AFF01FFFFA0FF00FF0000FF00FF3FFFFF00FFFC00FF";
    attribute INIT_1B of inst : label is "0000FFFF0000FFFF0000FFFF0000FFFFFFFF0000FFFF0000FFFFFF00FFFF00FF";
    attribute INIT_1C of inst : label is "000000FF0000FF00FFFF0000FFFF000000003FFF0000FFFC0AFF0000FFA00000";
    attribute INIT_1D of inst : label is "00FF0000FF000000000000FF0000FF00002F0000F800000000FF00FFFF00FF00";
    attribute INIT_1E of inst : label is "000000FF0000FF0001FFFFFFFF40FFFFFFFF00FFFFFFFF000000FFFF0000FFFF";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000FFFF00FFFFFFFF00002F0000F8000000";
    attribute INIT_20 of inst : label is "002F003F0010000AFE00FF000100A80000F700D7004000BECC003C0004007800";
    attribute INIT_21 of inst : label is "0FFF2FFF001F00AAFFF0FFF8FFD0000037FF01F700016A00F800FFE0F3FC0000";
    attribute INIT_22 of inst : label is "0000000000000000000000008000000003FF0FFF01510000F7C0FFF095000000";
    attribute INIT_23 of inst : label is "3FFF3FFF00000000FFFCFFFC00000000000303FF000100000000FF0000000000";
    attribute INIT_24 of inst : label is "3FFF1F0F01FF0A02F6FCC3F4FF4080A03FFF1F0F01FF2028F6FCC3F4FF402008";
    attribute INIT_25 of inst : label is "00FF000500000A80FF002CA0000002A00FFF000500002A00F8002CA000002A00";
    attribute INIT_26 of inst : label is "000000000000AAAA000000000000AAA0000000000000AAAA054000000000AAA0";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "3FFF07FF00030A00FFF0FF40000002803FFF07FF00030080FFF0FF4000000800";
    attribute INIT_2F of inst : label is "58D50C8300000000262633330000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "3FFF1FC301FF0A02FFFCF0F4FF4080A03FFF1FC301FF2028FFFCF0F4FF402808";
    attribute INIT_31 of inst : label is "3FFF1C0301FF0A02FFFCC034FF4080A03FFF1C0301FF2028FFFCC034FF402808";
    attribute INIT_32 of inst : label is "3FFF1F0F01FF0A02FFFCC3F4FF4080A03FFF1F0F01FF2028FFFCC3F4FF402808";
    attribute INIT_33 of inst : label is "3FFF1D0701FF0A02FFFCD074FF4080A03FFF1D0701FF2028FFFCD074FF402808";
    attribute INIT_34 of inst : label is "00C206C30000000058960CC3000000001D5220330000000058960CC300000000";
    attribute INIT_35 of inst : label is "C962CC230000000058960CC300000000256230330000000058960CC300000000";
    attribute INIT_36 of inst : label is "00003FE007FF000000002FF0FF4000000FFF3FE007FF000040000000E0000000";
    attribute INIT_37 of inst : label is "0FE03FFE07FF00002FC0FFF0FF4000000FFF3FFE07FF0000FFC08000FF400000";
    attribute INIT_38 of inst : label is "000000000000000000000000000000000FFF3FFF07FF0000FFC0FFF0FF400000";
    attribute INIT_39 of inst : label is "3FFF1D0701AF2028FFF0D074FA402AA83FFF1F5F000B2028FFF0F5F4E0002AA8";
    attribute INIT_3A of inst : label is "00A8BFFD10000000A800FFF80010000002BF3FF414000000FA007FF000500000";
    attribute INIT_3B of inst : label is "0AA0FF55000000002A8057FC0000000000A8FFF500000000A8007FFC00000000";
    attribute INIT_3C of inst : label is "BFFE000500000000FFF84000000000002BFE005500000000FFA0540000000000";
    attribute INIT_3D of inst : label is "007F000100000000F40000000000000017FF000100000000FF50000000000000";
    attribute INIT_3E of inst : label is "00030001000000000000000000000000000F000100000000C000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000400240000000000900080000000000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "155501E001543EAD1554000F00543D7D055502AD055407E8014003C001503C0F";
    attribute INIT_01 of inst : label is "15553EA815553EA815503C0F01543C0015543EAD01503D5F05540AAF05501AF5";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0F3C00000F3C000000000F0000000000000500AFFFC0E800000001FF0000FD00";
    attribute INIT_05 of inst : label is "00000000D000F00007FF0F007FFFF000FFD0F0F0D0FFF0F003FF0FAAFFFDF00F";
    attribute INIT_06 of inst : label is "3EAF03C007E83C0F3EA8140F01FC2ABE0ABE140F1EAD1F8007C003C006B42F0E";
    attribute INIT_07 of inst : label is "C000C000EAAAC00000030003AAAB000300000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D2F3EAA3C003EAA3C003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F2BE803C03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "000040000000C02A0000EA001AA4C94300FC02002ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "003F00000000003FFFFF00000000FF503FFF000000003FF40000000000000000";
    attribute INIT_0D of inst : label is "000000000000000001FF00000000000003FF0000000003FFFFFF00000000D400";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "00060001706930C391A4330CEAC60C0CEA8640CCAB8640CC0706030C00000000";
    attribute INIT_11 of inst : label is "00000000900030001A4630CCA8690CC3000E0004B8690CC3000A0004A46980C3";
    attribute INIT_12 of inst : label is "003F0000FF00C0000000003F0000FF0000390036B30073000000003E0000E700";
    attribute INIT_13 of inst : label is "0FFF0BFFFFF02A8000001FFF5500FFFC1BFF3FFAFF8000000000001B0545FFF8";
    attribute INIT_14 of inst : label is "003800033800800000050383580083800FFF00BEFCF0FE0000000FFF0000FFD0";
    attribute INIT_15 of inst : label is "3FFF0AFFFFFCFFA0000005F00000075000BB0003B80000000000001F0000D000";
    attribute INIT_16 of inst : label is "00000000000000003E2C000038BC00007050FFFC0FC13FFF0000F5000000005F";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000555500005555000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "FF00FFFF00FFFFFFFF003FFF00FFFFFCFF00FF0000FF00FF05FFFF80FF5002FF";
    attribute INIT_1B of inst : label is "0000FFFF0000FFFF0000FFFF0000FFFFFFFF0000FFFF0000FFFFFF80FFFF02FF";
    attribute INIT_1C of inst : label is "0000001F0000F400FFFF0000FFFF0000000005FF0000FF503FFF0000FFFC0000";
    attribute INIT_1D of inst : label is "00FF0000FF000000000000FF0000FF0000FF0000FF00000000FF00FFFF00FF00";
    attribute INIT_1E of inst : label is "0000001F0000F40000FFFFFFFF00FFFFFFFF02FFFFFFFF800000FFFF0000FFFF";
    attribute INIT_1F of inst : label is "00000000000000000000000000000000FFFF02FFFFFFFF8000FF0000FF000000";
    attribute INIT_20 of inst : label is "003F003F00000000FF00FF000000C00000E600FB000000D96C009C000000CC00";
    attribute INIT_21 of inst : label is "0FFF1FFF00000BFFFFF0FFFC55002A001BFF001B00003FFAFF80FFF805450000";
    attribute INIT_22 of inst : label is "003803830005000338008380580080000FFF0FFF000000BEFCF0FFD00000FE00";
    attribute INIT_23 of inst : label is "3FFF05F000000AFFFFFC07500000FFA000BB001F00000003B800D00000000000";
    attribute INIT_24 of inst : label is "3D7F082E00053FEF5E640BF05000F2FC3D7F082E00053EFE5E640BF05000B6BC";
    attribute INIT_25 of inst : label is "001F000000000FFFFF0014500000FFF001FF000000003FFFFE0014500000FF00";
    attribute INIT_26 of inst : label is "0000000000001F550000000000005FF40000000000001FD7000000000000FFF4";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "1FFF001700002FFAFFD050000000BFE01FFF001700002FEAFFD050000000AFE0";
    attribute INIT_2F of inst : label is "A418501400000000333304040000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "3FF50FE000053FEFFD7CB8205000FBFC3FF50FE000053EFEFD7CB8205000BFBC";
    attribute INIT_31 of inst : label is "3DF70FAF00053FEFDF7CFAF05000FBFC3DF70FAF00053EFEDF7CFAF05000BFBC";
    attribute INIT_32 of inst : label is "3D7F082E00053FEF5FFC0BF05000FBFC3D7F082E00053EFE5FFC0BF05000BFBC";
    attribute INIT_33 of inst : label is "3FFF0CA300053FEFFFFCCA305000FBFC3FFF0CA300053EFEFFFCCA305000BFBC";
    attribute INIT_34 of inst : label is "75D30040000000000CC350140000000001830540000000000CC3501400000000";
    attribute INIT_35 of inst : label is "CE934140000000000CC35014000000001A930540000000000CC3501400000000";
    attribute INIT_36 of inst : label is "3E001FFE0015000002F0FFD0500000003FF41FFE001502BF000000005000F000";
    attribute INIT_37 of inst : label is "3FF81FFF00150280BFF0FFD050000A003FFF1FFF001502BFD400FE805000FA00";
    attribute INIT_38 of inst : label is "000000000000000000000000000000003FFF1FFF001502BFFFF0FFD05000FA00";
    attribute INIT_39 of inst : label is "3FFF0C0300053EFEFFF0C0305000BFD43FFF0C0300053EFEFFF0C0305000BFD4";
    attribute INIT_3A of inst : label is "2FFFFF4000000000FFE007FC000000000FFF3F4000000000FFC007F000000000";
    attribute INIT_3B of inst : label is "BFFF000000000000FFF80000000000002FFF540000000000FFE0005400000000";
    attribute INIT_3C of inst : label is "15FF0000000002A0FD50000000002A00FFFF000000000000FFFC000000000000";
    attribute INIT_3D of inst : label is "001F0000000002FED00000000000FE00005F000000002FF8D40000000000BFE0";
    attribute INIT_3E of inst : label is "00030000000000030000000000000000000700000000002E400000000000E000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000005000024000002180280610000009000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
