library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_PROG_ROM_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_PROG_ROM_3 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FD",X"07",X"FE",X"06",X"FB",X"07",X"FC",X"3C",X"45",X"BC",X"45",X"5E",X"46",X"B4",X"46",X"00",
		X"10",X"80",X"AA",X"00",X"32",X"10",X"00",X"BF",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",X"0F",
		X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"A2",X"57",X"91",X"27",X"BD",X"A3",X"57",
		X"C8",X"91",X"27",X"20",X"38",X"78",X"28",X"60",X"98",X"38",X"65",X"27",X"85",X"27",X"90",X"02",
		X"E6",X"28",X"60",X"A5",X"1A",X"C9",X"80",X"90",X"11",X"49",X"FF",X"85",X"1A",X"A5",X"19",X"49",
		X"FF",X"69",X"00",X"85",X"19",X"90",X"02",X"E6",X"1A",X"38",X"26",X"37",X"A5",X"1C",X"C9",X"80",
		X"90",X"11",X"49",X"FF",X"85",X"1C",X"A5",X"1B",X"49",X"FF",X"69",X"00",X"85",X"1B",X"90",X"02",
		X"E6",X"1C",X"38",X"26",X"37",X"A5",X"19",X"C5",X"1B",X"A5",X"1A",X"E5",X"1C",X"A2",X"00",X"B0",
		X"02",X"A2",X"02",X"B5",X"1A",X"A0",X"09",X"C9",X"02",X"B0",X"09",X"88",X"16",X"19",X"F0",X"03",
		X"2A",X"10",X"F4",X"2A",X"95",X"1A",X"98",X"0A",X"66",X"37",X"2A",X"66",X"37",X"2A",X"0A",X"85",
		X"37",X"8A",X"49",X"02",X"AA",X"C0",X"09",X"B0",X"07",X"C8",X"16",X"19",X"36",X"1A",X"10",X"F5",
		X"A0",X"00",X"A5",X"1B",X"91",X"27",X"A5",X"37",X"29",X"FC",X"05",X"1C",X"C8",X"91",X"27",X"A5",
		X"19",X"C8",X"91",X"27",X"A5",X"37",X"29",X"02",X"0A",X"05",X"8F",X"05",X"1A",X"C8",X"91",X"27",
		X"4C",X"38",X"78",X"A2",X"02",X"BD",X"01",X"24",X"0A",X"B5",X"B7",X"29",X"1F",X"B0",X"37",X"F0",
		X"10",X"C9",X"1B",X"B0",X"0A",X"A8",X"A5",X"BA",X"29",X"07",X"C9",X"07",X"98",X"90",X"02",X"E9",
		X"01",X"95",X"B7",X"AD",X"00",X"20",X"29",X"04",X"D0",X"04",X"A9",X"F0",X"85",X"B4",X"A5",X"B4",
		X"F0",X"08",X"C6",X"B4",X"A9",X"00",X"95",X"B7",X"95",X"B3",X"18",X"B5",X"B3",X"F0",X"23",X"D6",
		X"B3",X"D0",X"1F",X"38",X"B0",X"1C",X"C9",X"1B",X"B0",X"09",X"B5",X"B7",X"69",X"20",X"90",X"D1",
		X"F0",X"01",X"18",X"A9",X"1F",X"B0",X"CA",X"95",X"B7",X"B5",X"B3",X"F0",X"01",X"38",X"A9",X"78",
		X"95",X"B3",X"90",X"04",X"F6",X"B6",X"E6",X"B2",X"CA",X"CA",X"10",X"99",X"E6",X"BA",X"A5",X"BA",
		X"4A",X"A5",X"B2",X"B0",X"0C",X"F0",X"0A",X"C9",X"10",X"B0",X"02",X"69",X"FF",X"69",X"EF",X"85",
		X"B2",X"0A",X"60",X"25",X"89",X"86",X"3C",X"05",X"3C",X"8D",X"00",X"3C",X"85",X"89",X"60",X"25",
		X"88",X"86",X"3C",X"05",X"3C",X"8D",X"00",X"32",X"85",X"88",X"60",X"AD",X"03",X"28",X"29",X"03",
		X"AA",X"BD",X"9B",X"79",X"85",X"99",X"A2",X"00",X"EE",X"00",X"58",X"F0",X"06",X"AD",X"02",X"28",
		X"29",X"03",X"AA",X"86",X"21",X"38",X"AD",X"01",X"28",X"2A",X"2A",X"2D",X"00",X"28",X"29",X"0F",
		X"69",X"00",X"C9",X"09",X"90",X"02",X"A9",X"00",X"85",X"98",X"60",X"01",X"04",X"05",X"06",X"A2",
		X"0C",X"A5",X"98",X"18",X"69",X"18",X"20",X"34",X"7A",X"A9",X"17",X"20",X"4F",X"7A",X"A9",X"05",
		X"20",X"4F",X"7A",X"A5",X"86",X"29",X"20",X"F0",X"07",X"A2",X"00",X"A9",X"04",X"4C",X"34",X"7A",
		X"60",X"00",X"84",X"37",X"A0",X"0F",X"86",X"38",X"A9",X"00",X"85",X"92",X"85",X"93",X"85",X"94",
		X"F8",X"06",X"37",X"26",X"38",X"A5",X"92",X"65",X"92",X"85",X"92",X"A5",X"93",X"65",X"93",X"85",
		X"93",X"A5",X"94",X"65",X"94",X"85",X"94",X"88",X"10",X"E7",X"A4",X"94",X"A6",X"93",X"A5",X"92",
		X"D8",X"60",X"86",X"2C",X"84",X"2B",X"A9",X"00",X"4A",X"A8",X"B1",X"2B",X"85",X"39",X"29",X"7F",
		X"AA",X"98",X"0A",X"A8",X"BD",X"A2",X"57",X"91",X"27",X"C8",X"BD",X"A3",X"57",X"91",X"27",X"C8",
		X"98",X"24",X"39",X"10",X"E3",X"18",X"65",X"27",X"85",X"27",X"90",X"02",X"E6",X"28",X"98",X"4A",
		X"65",X"2B",X"85",X"2B",X"90",X"02",X"E6",X"2C",X"60",X"A9",X"17",X"20",X"4F",X"7A",X"A9",X"03",
		X"D0",X"1D",X"A9",X"80",X"48",X"8A",X"18",X"69",X"0C",X"A8",X"A9",X"55",X"69",X"00",X"A6",X"27",
		X"86",X"2F",X"A6",X"28",X"86",X"30",X"20",X"CD",X"7E",X"20",X"10",X"7F",X"68",X"30",X"58",X"C9",
		X"18",X"90",X"03",X"0A",X"D0",X"48",X"48",X"A6",X"21",X"F0",X"10",X"CA",X"7D",X"A1",X"5F",X"AA",
		X"BD",X"A4",X"5F",X"A2",X"00",X"0A",X"90",X"0F",X"CA",X"B0",X"0C",X"E9",X"08",X"C9",X"0C",X"B0",
		X"13",X"AA",X"BD",X"6D",X"69",X"A2",X"00",X"18",X"A0",X"02",X"71",X"2F",X"91",X"2F",X"8A",X"C8",
		X"71",X"2F",X"91",X"2F",X"68",X"0A",X"C9",X"30",X"B0",X"14",X"A6",X"21",X"F0",X"10",X"CA",X"18",
		X"7D",X"00",X"58",X"AA",X"BC",X"04",X"58",X"BD",X"05",X"58",X"AA",X"4C",X"F2",X"79",X"AA",X"BC",
		X"2B",X"69",X"BD",X"2C",X"69",X"D0",X"F3",X"60",X"48",X"8A",X"48",X"98",X"48",X"D8",X"AD",X"00",
		X"2C",X"38",X"E5",X"83",X"B0",X"04",X"C6",X"83",X"A9",X"00",X"C5",X"84",X"90",X"04",X"E6",X"84",
		X"A5",X"84",X"AA",X"38",X"E5",X"82",X"90",X"0A",X"4A",X"4A",X"F0",X"0A",X"86",X"82",X"E6",X"85",
		X"D0",X"04",X"69",X"03",X"30",X"F6",X"E6",X"74",X"A5",X"73",X"C9",X"03",X"B0",X"0D",X"8D",X"00",
		X"34",X"A5",X"00",X"45",X"C1",X"45",X"C2",X"C9",X"85",X"F0",X"03",X"4C",X"EB",X"7A",X"20",X"D3",
		X"78",X"90",X"06",X"A2",X"20",X"A9",X"FF",X"D0",X"04",X"A9",X"DF",X"A2",X"00",X"20",X"5F",X"79",
		X"24",X"22",X"50",X"2F",X"C6",X"87",X"D0",X"2B",X"A9",X"FA",X"85",X"87",X"E6",X"8D",X"F8",X"18",
		X"A2",X"00",X"A0",X"02",X"A9",X"08",X"75",X"9E",X"95",X"9E",X"A9",X"00",X"E8",X"88",X"10",X"F6",
		X"A5",X"9C",X"18",X"69",X"01",X"C9",X"60",X"90",X"02",X"A9",X"00",X"85",X"9C",X"A5",X"9D",X"69",
		X"00",X"85",X"9D",X"D8",X"A5",X"22",X"D0",X"0E",X"A5",X"74",X"A2",X"1F",X"4A",X"90",X"02",X"A2",
		X"10",X"A9",X"00",X"20",X"5F",X"79",X"C6",X"8A",X"D0",X"06",X"A9",X"06",X"85",X"8A",X"E6",X"73",
		X"68",X"A8",X"68",X"AA",X"68",X"40",X"00",X"A0",X"02",X"38",X"08",X"88",X"84",X"38",X"18",X"65",
		X"38",X"28",X"AA",X"08",X"86",X"37",X"B5",X"00",X"4A",X"4A",X"4A",X"4A",X"28",X"20",X"18",X"78",
		X"A5",X"38",X"D0",X"01",X"18",X"A6",X"37",X"B5",X"00",X"20",X"18",X"78",X"A6",X"37",X"CA",X"C6",
		X"38",X"10",X"E0",X"60",X"A2",X"FF",X"9A",X"D8",X"A9",X"00",X"8D",X"00",X"3C",X"AA",X"95",X"00",
		X"E8",X"D0",X"FB",X"AD",X"00",X"20",X"4A",X"4A",X"B0",X"03",X"4C",X"B9",X"7B",X"A9",X"85",X"85",
		X"00",X"85",X"C1",X"85",X"C2",X"A9",X"FF",X"85",X"83",X"A9",X"06",X"85",X"8A",X"A9",X"02",X"85",
		X"9A",X"85",X"9B",X"8D",X"00",X"34",X"4C",X"01",X"60",X"A2",X"11",X"9A",X"8A",X"85",X"00",X"A0",
		X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"D0",X"23",X"E8",X"D0",X"F7",X"BA",X"8A",X"8D",X"00",
		X"34",X"C8",X"D9",X"00",X"00",X"D0",X"12",X"A2",X"00",X"96",X"00",X"C8",X"D0",X"05",X"0A",X"A2",
		X"00",X"B0",X"0A",X"AA",X"9A",X"96",X"00",X"D0",X"D8",X"59",X"00",X"00",X"AA",X"8A",X"A0",X"10",
		X"29",X"0F",X"F0",X"02",X"A0",X"20",X"8A",X"A2",X"10",X"29",X"F0",X"F0",X"02",X"A2",X"20",X"98",
		X"9A",X"AA",X"8E",X"00",X"3C",X"A0",X"0C",X"A2",X"64",X"2C",X"00",X"20",X"70",X"FB",X"2C",X"00",
		X"20",X"50",X"FB",X"8D",X"00",X"34",X"CA",X"D0",X"F0",X"C0",X"05",X"D0",X"03",X"8E",X"00",X"3C",
		X"88",X"D0",X"E4",X"A8",X"30",X"05",X"09",X"80",X"BA",X"10",X"D7",X"C9",X"90",X"D0",X"05",X"BA",
		X"E0",X"10",X"F0",X"06",X"8D",X"00",X"34",X"4C",X"34",X"7C",X"A2",X"FF",X"9A",X"20",X"59",X"7E",
		X"A8",X"91",X"27",X"C8",X"D0",X"FB",X"E6",X"28",X"A6",X"28",X"E0",X"48",X"90",X"F3",X"20",X"59",
		X"7E",X"A9",X"11",X"85",X"37",X"84",X"BC",X"91",X"27",X"98",X"AA",X"C8",X"F0",X"06",X"B1",X"27",
		X"D0",X"2B",X"F0",X"F7",X"8A",X"A8",X"A5",X"37",X"8D",X"00",X"34",X"D1",X"27",X"D0",X"1C",X"A9",
		X"00",X"91",X"27",X"A5",X"37",X"C8",X"D0",X"03",X"0A",X"B0",X"06",X"85",X"37",X"91",X"27",X"D0",
		X"D8",X"E6",X"28",X"A5",X"28",X"C9",X"48",X"90",X"C8",X"B0",X"1E",X"51",X"27",X"A2",X"00",X"48",
		X"29",X"F0",X"F0",X"02",X"A2",X"02",X"68",X"29",X"0F",X"F0",X"01",X"E8",X"8A",X"A6",X"28",X"E0",
		X"44",X"90",X"02",X"0A",X"0A",X"05",X"BC",X"85",X"BC",X"A5",X"BC",X"8D",X"00",X"32",X"A9",X"03",
		X"85",X"56",X"18",X"A9",X"10",X"66",X"BC",X"08",X"90",X"01",X"0A",X"8D",X"00",X"3C",X"A0",X"50",
		X"20",X"7F",X"7E",X"8E",X"00",X"3C",X"A0",X"28",X"20",X"7F",X"7E",X"28",X"C6",X"56",X"10",X"E3",
		X"66",X"BC",X"8D",X"00",X"34",X"D0",X"FB",X"A9",X"48",X"85",X"2C",X"20",X"59",X"7E",X"85",X"2B",
		X"85",X"BC",X"85",X"BB",X"20",X"2D",X"7F",X"A9",X"12",X"20",X"62",X"7E",X"A2",X"37",X"8A",X"0A",
		X"A0",X"00",X"8D",X"00",X"34",X"51",X"2B",X"C8",X"D0",X"FB",X"A8",X"8A",X"29",X"03",X"C9",X"01",
		X"98",X"B0",X"2E",X"F0",X"2B",X"85",X"BC",X"86",X"39",X"A9",X"34",X"38",X"E5",X"39",X"4A",X"85",
		X"3A",X"38",X"E9",X"04",X"C9",X"04",X"B0",X"02",X"C6",X"BB",X"A5",X"BC",X"29",X"0F",X"F0",X"03",
		X"20",X"17",X"7F",X"A5",X"BC",X"29",X"F0",X"F0",X"05",X"E6",X"3A",X"20",X"17",X"7F",X"A6",X"39",
		X"8A",X"E6",X"2C",X"CA",X"10",X"BA",X"A6",X"BC",X"F0",X"16",X"24",X"BB",X"10",X"1B",X"A9",X"40",
		X"85",X"27",X"A9",X"18",X"85",X"27",X"A9",X"22",X"A2",X"0E",X"20",X"64",X"7E",X"4C",X"59",X"7D",
		X"AE",X"7F",X"7F",X"AC",X"7E",X"7F",X"20",X"F2",X"79",X"A9",X"00",X"85",X"56",X"85",X"39",X"85",
		X"89",X"A9",X"11",X"8D",X"00",X"32",X"A5",X"28",X"85",X"2A",X"A5",X"27",X"85",X"29",X"A2",X"07",
		X"BD",X"00",X"24",X"0A",X"26",X"BD",X"CA",X"10",X"F7",X"AD",X"00",X"20",X"29",X"04",X"85",X"BE",
		X"A2",X"00",X"A5",X"BF",X"45",X"BD",X"D0",X"06",X"A5",X"C0",X"45",X"BE",X"F0",X"02",X"A2",X"30",
		X"A9",X"0F",X"20",X"53",X"79",X"A5",X"BD",X"85",X"BF",X"A5",X"BE",X"85",X"C0",X"A5",X"29",X"85",
		X"27",X"A5",X"2A",X"85",X"28",X"24",X"BB",X"30",X"27",X"A9",X"1A",X"20",X"62",X"7E",X"A0",X"01",
		X"AD",X"00",X"2C",X"18",X"65",X"82",X"6A",X"85",X"82",X"A9",X"82",X"20",X"59",X"7B",X"20",X"9F",
		X"79",X"A9",X"3A",X"20",X"62",X"7E",X"20",X"6B",X"79",X"A9",X"99",X"A0",X"01",X"20",X"59",X"7B",
		X"20",X"71",X"7E",X"E6",X"56",X"A5",X"56",X"C9",X"20",X"90",X"1C",X"A6",X"3A",X"E8",X"E0",X"05",
		X"90",X"02",X"A2",X"00",X"86",X"3A",X"BD",X"80",X"7F",X"8D",X"00",X"32",X"BD",X"85",X"7F",X"AA",
		X"A9",X"30",X"20",X"53",X"79",X"84",X"56",X"20",X"95",X"7E",X"B0",X"03",X"4C",X"6E",X"7D",X"A2",
		X"00",X"8E",X"00",X"3C",X"86",X"BB",X"20",X"59",X"7E",X"A4",X"BB",X"C0",X"03",X"D0",X"23",X"A9",
		X"30",X"20",X"62",X"7E",X"A9",X"FB",X"A0",X"00",X"91",X"27",X"E6",X"27",X"48",X"A9",X"F8",X"91",
		X"27",X"E6",X"27",X"A9",X"38",X"A2",X"02",X"20",X"64",X"7E",X"68",X"38",X"E9",X"10",X"B0",X"E6",
		X"90",X"12",X"BE",X"F4",X"7F",X"98",X"0A",X"A8",X"B9",X"EF",X"7F",X"48",X"B9",X"EE",X"7F",X"A8",
		X"68",X"20",X"A6",X"7E",X"20",X"71",X"7E",X"20",X"7A",X"7E",X"20",X"95",X"7E",X"90",X"F8",X"A6",
		X"BB",X"E8",X"E0",X"04",X"90",X"AE",X"4C",X"9D",X"7B",X"A9",X"40",X"85",X"28",X"A9",X"00",X"85",
		X"27",X"60",X"A2",X"08",X"18",X"6D",X"7C",X"7F",X"A8",X"AD",X"7D",X"7F",X"69",X"00",X"4C",X"A6",
		X"7E",X"A9",X"4B",X"A0",X"DE",X"A2",X"06",X"20",X"A6",X"7E",X"8D",X"00",X"30",X"A0",X"03",X"8D",
		X"00",X"34",X"A2",X"14",X"2C",X"00",X"20",X"70",X"FB",X"2C",X"00",X"20",X"50",X"FB",X"CA",X"D0",
		X"F3",X"88",X"D0",X"EB",X"60",X"2C",X"00",X"20",X"30",X"03",X"06",X"26",X"60",X"A9",X"20",X"85",
		X"26",X"18",X"90",X"F8",X"A2",X"08",X"85",X"65",X"84",X"64",X"8A",X"A8",X"88",X"B1",X"64",X"91",
		X"27",X"88",X"10",X"F9",X"8A",X"18",X"65",X"27",X"85",X"27",X"90",X"02",X"E6",X"28",X"8A",X"18",
		X"65",X"64",X"85",X"64",X"90",X"02",X"E6",X"65",X"60",X"A2",X"02",X"D0",X"D9",X"A2",X"04",X"D0",
		X"D5",X"A2",X"04",X"D0",X"D5",X"18",X"65",X"8B",X"A8",X"8A",X"69",X"00",X"A2",X"00",X"86",X"3D",
		X"A2",X"0F",X"86",X"3E",X"85",X"65",X"84",X"64",X"A0",X"00",X"B1",X"64",X"38",X"E5",X"53",X"91",
		X"27",X"C8",X"B1",X"64",X"E5",X"54",X"29",X"0F",X"09",X"A0",X"91",X"27",X"C8",X"B1",X"64",X"38",
		X"E5",X"51",X"91",X"27",X"C8",X"B1",X"64",X"E5",X"3D",X"25",X"3E",X"91",X"27",X"20",X"38",X"78",
		X"A9",X"55",X"A0",X"AE",X"4C",X"CD",X"7E",X"A2",X"00",X"A4",X"3A",X"20",X"C2",X"79",X"A9",X"92",
		X"38",X"A0",X"01",X"20",X"5A",X"7B",X"A9",X"10",X"A2",X"02",X"4C",X"64",X"7E",X"A9",X"00",X"A2",
		X"10",X"4C",X"64",X"7E",X"00",X"A0",X"00",X"00",X"00",X"90",X"00",X"00",X"FF",X"A2",X"FF",X"03",
		X"00",X"90",X"00",X"00",X"0B",X"F0",X"58",X"A2",X"10",X"00",X"00",X"70",X"00",X"00",X"80",X"A1",
		X"00",X"02",X"00",X"70",X"00",X"00",X"CB",X"F8",X"C8",X"FF",X"CF",X"F8",X"C8",X"FB",X"CB",X"FF",
		X"0F",X"F8",X"CB",X"FB",X"90",X"A1",X"00",X"02",X"00",X"90",X"00",X"00",X"0F",X"FD",X"F4",X"A1",
		X"76",X"01",X"00",X"70",X"00",X"00",X"38",X"32",X"2E",X"00",X"32",X"AA",X"34",X"7F",X"76",X"7F",
		X"11",X"12",X"14",X"18",X"00",X"01",X"03",X"07",X"0F",X"00",X"80",X"A1",X"00",X"02",X"00",X"90",
		X"00",X"00",X"20",X"73",X"20",X"C3",X"07",X"E0",X"00",X"A0",X"00",X"00",X"00",X"90",X"00",X"00",
		X"FF",X"92",X"FF",X"C2",X"FC",X"77",X"FC",X"C3",X"FE",X"87",X"FE",X"C7",X"FE",X"83",X"FE",X"C7",
		X"FC",X"73",X"FC",X"C3",X"FF",X"96",X"FF",X"C2",X"FF",X"92",X"01",X"00",X"FF",X"96",X"FF",X"C6",
		X"FC",X"73",X"FC",X"C7",X"FE",X"83",X"FE",X"C3",X"FE",X"87",X"FE",X"C3",X"FC",X"77",X"FC",X"C7",
		X"FF",X"92",X"FF",X"C6",X"80",X"A1",X"00",X"02",X"00",X"90",X"00",X"00",X"06",X"C0",X"00",X"B0",
		X"08",X"C0",X"00",X"D0",X"0A",X"C0",X"00",X"D0",X"CB",X"FB",X"CF",X"FB",X"00",X"D0",X"8A",X"7F",
		X"98",X"7F",X"D4",X"7F",X"0E",X"3C",X"1A",X"00",X"57",X"00",X"A8",X"7A",X"84",X"7B",X"84",X"7B");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
