-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "98384A5BC6C110B665C263A0A1A90ED87E2716DDF425B396BF50AFD6F4261059";
    attribute INIT_01 of inst : label is "4B25CDB36DB9E2717480E3339E2102802534016317213FF6C8B2934B6DD3C249";
    attribute INIT_02 of inst : label is "036DCCCD2D11BB37C034CE7D69DAF52FB72DF735D034CDF9F24CC47D5D573572";
    attribute INIT_03 of inst : label is "CB7D3C64CD37FBB9B729603C9AEB588832CF67314D4FABFDFF73CF6C4B35145A";
    attribute INIT_04 of inst : label is "3708DD63126161358C8E831988AD7018C4E74D343FDDC0C87293A4F37F6F90B3";
    attribute INIT_05 of inst : label is "B22B0BCB7CE827043FD603C62E7A0292737D08CFE9D3CC8B98892E733A9CA0E3";
    attribute INIT_06 of inst : label is "9E398CA69999898626AAEABFC10C0A6A7495ED694555357AAF68D65811844313";
    attribute INIT_07 of inst : label is "5F6D6D53180AFBAF57DFF57FEBEAEF9800E270E7420CDA2FD9996E6599F9B9F9";
    attribute INIT_08 of inst : label is "73954C33A0AFCFC76E750105A0C886245003CB91E62EF37E3C13BCF89EBF37F0";
    attribute INIT_09 of inst : label is "1E7140B4178B3A2E313123264BBA66AE02C3777137EC71F9D49B347114F9FD63";
    attribute INIT_0A of inst : label is "7FDCEF9DEF68FB11E29A73FBE64DB2DBBC06E119A0E6B19845F4477459BDF21B";
    attribute INIT_0B of inst : label is "05B9B045DF98791C62188721DE450024219DB9FFAE6778D7FF1E3E3FCFCEFFDA";
    attribute INIT_0C of inst : label is "331C3330F62A252405030F9D8C9F608B4E8965CCDE528F2DE2F4EE272F775CA0";
    attribute INIT_0D of inst : label is "1C8D363719E6639E053E6D33AE266B6E4D9A36A4B6FE7DF388D35E0497609584";
    attribute INIT_0E of inst : label is "8A8CC0884674BB46CAB48C89F7961E9A3ED0C44912314E2D8D17BE2D8DCDD597";
    attribute INIT_0F of inst : label is "91CF0F9987F604AB1434D8CD5F998807A8CC0B270DF6223AC725633B0C1AED92";
    attribute INIT_10 of inst : label is "3636E6463A7C665CBC21A5E5679BAE4253302FCF4BADF7A122302F6CB23AA960";
    attribute INIT_11 of inst : label is "FE88F306FBF248C734FC6CF2EFC4EB2049C8FDFF0A19A94A1D24DDD9BB647340";
    attribute INIT_12 of inst : label is "33EE5B5FAE6E619A7D10D4D52322322234CC041741578DA13543B596D1792F24";
    attribute INIT_13 of inst : label is "303D779E864A6C9AF0FC221769A7AE9734D92D33093261BC0D074341BB558654";
    attribute INIT_14 of inst : label is "0D3DE4EAD969AF6C44519BA346859595AD07AF0C9288D2CA0B0B0F0FCACACACB";
    attribute INIT_15 of inst : label is "8478F1F7E78F22B83D50FC9D67632A636CD760D869FDA3F727D75CDEC9AD121D";
    attribute INIT_16 of inst : label is "DC1D5FDCE0B97CEE413535949CA7E4A3C6361C2234CB4D09E3D10DE2D9BE7820";
    attribute INIT_17 of inst : label is "821F4D515FF3CF55AE32E4D0DF5DF58DD787E7DDAE6ABDE2CF828CF3525C2D1D";
    attribute INIT_18 of inst : label is "6FFDCA4FFE50212AF02BF216E1AB4AF7FAFAFEB5F32DE23FB2F60088FB65F7A0";
    attribute INIT_19 of inst : label is "DB6CF7CF665B6F97CBFF3CB3F9C69FAAF77CF2B1F3DC5AAF364DE1C66CF0EFFB";
    attribute INIT_1A of inst : label is "FC8CDDD89B8297FBB4C1BCBD13E7B7E70CC837DCD004D23C72379CF6CF4F21F3";
    attribute INIT_1B of inst : label is "CFD529D95D6CFEFEF4A05B3C9DCBA74F6CCD06C8FB6FFD69F24A43CF077759EF";
    attribute INIT_1C of inst : label is "1810464D80A8ACE8145590150AB230A8BCD25208C7D6C9ADD74F82737FB53C1F";
    attribute INIT_1D of inst : label is "55850506A210B4AA1C425C5CA8A8A801559618407730F4F99D151D95022DC4E5";
    attribute INIT_1E of inst : label is "511C4105CF36DEDB000050407195FD4A550094B577939551505141415561F404";
    attribute INIT_1F of inst : label is "4F98CEDDBAC6584A4514542F679BD899712D53452D172C7551984551E646E4B5";
    attribute INIT_20 of inst : label is "ECB262F71AE501F73CF36F43B38C7E55017C69F29D8C502765F3F1CB7E7BDD68";
    attribute INIT_21 of inst : label is "98FF2320F18D43FD43CC27C55B60DFED20E51FFD679EA799953F3DDD3023326B";
    attribute INIT_22 of inst : label is "B0155005A93544F08DE6809E6E24948510037036B0D3FFC4F630277374ECE35D";
    attribute INIT_23 of inst : label is "F963796E95DDEFD3F5E35A6DB008DFE0CE5C88BF3F45D4738E415D722C30DDDB";
    attribute INIT_24 of inst : label is "090088005CD55244919DE7960194B2B0912358E121A37DD534D24D74FDFDD379";
    attribute INIT_25 of inst : label is "F7BCE3D6088E907E59BD3CF2F0A021CCC938F78D40CF1930D32FF6364C0F1A2C";
    attribute INIT_26 of inst : label is "D0986732CFAAD76F4FB3CB66CE5E7F4FFE95555A15555552EB2F9BF7D9DE7EEF";
    attribute INIT_27 of inst : label is "C771DC0F6207F5E67D9C83F23CE3F60F5D3234C3C4AA338CC6C4A1FF4C50E8C8";
    attribute INIT_28 of inst : label is "9C7027189FA1FFB02025DF011709A98E0C909C74FCBF754771CC1FC44FF87675";
    attribute INIT_29 of inst : label is "ACB866137EFEA3B364B0A498FEA717F7BF4D33A4D3BDF4B9C21C258751F72950";
    attribute INIT_2A of inst : label is "6E99C97DA3369F3C3992D2CDBCD26B0A66872AD3A754D5F75329DFD0DBC99D8B";
    attribute INIT_2B of inst : label is "9477131FA80D837C7734432BE1D6E2593754DD7DC16F14F4C894B90EC1B66DD9";
    attribute INIT_2C of inst : label is "B6DB2526D927BAED14F6DD2712EE204CC2676F0FED63DD6C2C20B13A62620BB3";
    attribute INIT_2D of inst : label is "DD8D2E3D878330EE090D9F6C97990CAE26018A5E109342F498242001F9F37924";
    attribute INIT_2E of inst : label is "CB3CF3C96EFC8FCBE44C3B766DB118749264F6CFF5771646A5348C455D71AFEB";
    attribute INIT_2F of inst : label is "3F0D438A9ED8BB2F7356E4E5229337D7CF53FB21241DF92535577CFD0D0547F2";
    attribute INIT_30 of inst : label is "2836358DA8CD21F92B17986FCEF3636BB50DF1333197689D6B5984366AABD28B";
    attribute INIT_31 of inst : label is "B6BBFD877B7B6F936CB793E0CB01BC6FBE43389BF6F7FCE0504D34C9CC1F3E77";
    attribute INIT_32 of inst : label is "B5DC4375A2C58CCF618DDCF51F162F9CACC8CFD27918D57B225918C44C955624";
    attribute INIT_33 of inst : label is "2EC810624F6DD037D575E3F373B75B3434CB51DF6F69DD8DB1F1F5BF45315DBC";
    attribute INIT_34 of inst : label is "DC04F575483CE8B981AD1C01619967DB0F831C5C54B5B4B1D484D5D4B4B962FC";
    attribute INIT_35 of inst : label is "5044551025B0E8310F5DC9E0868242BAE04C24DD2110DCAF036F10C3956BBA6F";
    attribute INIT_36 of inst : label is "171CCA73E76DA62D51441110261A027696CD5791BDB0F1F109111915A1B181B0";
    attribute INIT_37 of inst : label is "F157055F9BBEBB9B855A1578EEEEFF2B01531554D05511D574434424E6E1BD51";
    attribute INIT_38 of inst : label is "444505858ACCA0A7A1156445A0A2A2A1A84405FEB1C450D117152D4598F451F0";
    attribute INIT_39 of inst : label is "2F279C4FB8EE2CB255440C7008679E1B6EDFDDB482CDF5F555405555806431F4";
    attribute INIT_3A of inst : label is "43C53EA4FF2E2AB157515555AAAEABABC5551C71557035F55551557555555557";
    attribute INIT_3B of inst : label is "A586EE974BF15178134C35D4ADCBFAB70D750850F4B4BC9747D2383493EB25BF";
    attribute INIT_3C of inst : label is "23E36DD5BAA8838C2D84DCC238CEB07103D90E086CA40441052CB3DD75B6D1C0";
    attribute INIT_3D of inst : label is "034D2503A1A3A0609345A8A7AB44E11765C186A9E694F0F00505851F70F07A70";
    attribute INIT_3E of inst : label is "B2585646DCFA50EB3BFDE3EDE9F3F02A55F95555D5595F9FF7155553907B15C5";
    attribute INIT_3F of inst : label is "556FCE658CB6B632E62274D970B8A234B1678DCBEAF70A74F55A230B09267775";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "526365C7DDC7C424CC68CDE87531538986C8C815F228BDDCC7F9053068280353";
    attribute INIT_01 of inst : label is "F519364DB0E6AE1408992DC909FCD542CA4283B5B3B3B8EA322CB931274DDC22";
    attribute INIT_02 of inst : label is "DAD2155314B968CAC18E14AD0C2AB912CC934CDE700E379AB8E3333063901B88";
    attribute INIT_03 of inst : label is "04D052A232C89CF70C9FDFC22585B190CC10DCD2D390D4214CC90042B0C86E21";
    attribute INIT_04 of inst : label is "0D4A32E90778B468B7316BD944F9786466DD15C573C2ABA2184D160564E4AC1D";
    attribute INIT_05 of inst : label is "C8B0B0654993B452AD64DF66BFE6ECFFFF02E7134A4296812F9218BFB1862B42";
    attribute INIT_06 of inst : label is "F9BFFA141319130B4E00A008448C525AFB5FB342495B375FD7BF68CC5A726C1C";
    attribute INIT_07 of inst : label is "FDD7FE6822FA8232FEB117C18CEA0882DD1BA7AFB33140A63BE64D9D2787C5C5";
    attribute INIT_08 of inst : label is "8C0BA3DD55F7B3B1C5DFA7BFF7F728496D6D343A60DA8833CF29C30FF8F0FE5E";
    attribute INIT_09 of inst : label is "D1DBB7C95E6ECD99A5956F95B0F5B99DD937EC07BA93A3D01CA39F00F91AC35D";
    attribute INIT_0A of inst : label is "FF7F3F7FA9F6F2BB5F57FDE56EB2FBEE5AB56AF78FF63FFAF64BDDCBD73F2929";
    attribute INIT_0B of inst : label is "37FB8DDDB778DEF7B5EDFB76B3ADF8FB7CBF57C6DD5F17FD3DBDD7DE1ED5E79F";
    attribute INIT_0C of inst : label is "276064C0C8EC3063625A7252B069CF0794F6DC13239DA0C63E8304D85E2DF706";
    attribute INIT_0D of inst : label is "F904B7CD5D0982202080E048C9190C19F2214B30005402292420019840B952FE";
    attribute INIT_0E of inst : label is "F1675A7FFEF3B8B2DD5623E761CE2BAAB75A54A672167030E34D45B0C3590364";
    attribute INIT_0F of inst : label is "766DD731BAFAFAEAF20024604FA9BA661635A58D93CDD8736195918D97D560F5";
    attribute INIT_10 of inst : label is "C95D20A4C8A513A40244A464760608B089C6C1C99BE3A4F839C6C1D4ACD1E056";
    attribute INIT_11 of inst : label is "18AA4DBA8F877C379503C24A9CDC9FD004D50781B3BCF73373153595B0E984E2";
    attribute INIT_12 of inst : label is "AF3191B6419AC02446F1773711001001A035D8DD3D69081880E4D9389A011059";
    attribute INIT_13 of inst : label is "8F85DF3D80548F24DE779C84104B2508953097D5635C18876EC1DFB08A766219";
    attribute INIT_14 of inst : label is "1603C48A96F4F88858577C1B1049F8AF17BD171DF64DF248F658B61A09060803";
    attribute INIT_15 of inst : label is "7D44051434E0D3F049782E0714B8E02E50708D37CED0BC6BC52C9E7EB0F2F052";
    attribute INIT_16 of inst : label is "2B805312425EBAA5B88C082E4078D0D0028101ED8F901BE25A00225B4450870A";
    attribute INIT_17 of inst : label is "28E121BA2D9FAAB978DD092F2D925933684C4D67D8B520959D796147E7EB2042";
    attribute INIT_18 of inst : label is "7AAD40B401741F608BDE0A002F2010A0CA8DAD8B5CD35AF5050A613DF4F628FF";
    attribute INIT_19 of inst : label is "24100D33B8A29861148CD249263161308D820C0CA8162ED0C4BF9828830E00AE";
    attribute INIT_1A of inst : label is "965F4753E9EDE724A5773271ECA8C93ABB455D667FB471E55E911A5C9DC5FF51";
    attribute INIT_1B of inst : label is "653E86753EBBC80E4E175D80CA2CE2F8174559456D15319C5E2E054537DDE664";
    attribute INIT_1C of inst : label is "87EBA5F8B5F0F5A5DEEF7FDFCDE7D38AFAFA487828069AC00F214D4C4A8C83C4";
    attribute INIT_1D of inst : label is "BF3F8BFDB01235F5E7BDAEA8EAEBF414BFB5E7ABF8FA1AFA0FA7AF0D7DF3DFEE";
    attribute INIT_1E of inst : label is "F4F779E7EBAEFEFBF3CF43F9BF83BFC2FFFB7FFF6D75BFFF657BF3F057DBFF7F";
    attribute INIT_1F of inst : label is "65267E63AACEABF2E79E7C1DEF8EFEACDFDBBDEFFB5DD7F7F4F4F7BFF34A5E7B";
    attribute INIT_20 of inst : label is "0040CD0855FA62E1F3094720CEBCB91274D4C1017FD3D3BDCD094F1B6442934B";
    attribute INIT_21 of inst : label is "7706CACAE3543DA5A4D0DD3A2EA621A5CB4A21A76C08AC83A0EF5E0929797CE0";
    attribute INIT_22 of inst : label is "AEFBEEBE906748FC6D2C43BFFBBE5392B001CEC8132434BA4007DC9CA2AA0917";
    attribute INIT_23 of inst : label is "2719CBA01A2889640831CF46C93302D320D3364C5392E1816A64134042EE36C8";
    attribute INIT_24 of inst : label is "575C72B15F43849BA6374F6674E6A5387D09F60D20B93396D6443305FA6AFD40";
    attribute INIT_25 of inst : label is "7D0F29A070F6C7312743DC453F39433B964BADF76ECFA76F78C01C796ECFB7AF";
    attribute INIT_26 of inst : label is "5D2F1AEB05BB59E2C449259B48BF7FAAD6FFFFF25F5F5F5AD4D4EF0CC2177DF3";
    attribute INIT_27 of inst : label is "A4A10A3C093095C2423A78C7FAAABA760EC1952C59DF40D25CEECE50458DAF61";
    attribute INIT_28 of inst : label is "0ACE82F7E85628545B4F6002C45AFA51F33E03E213C10AA0E9286C003082080B";
    attribute INIT_29 of inst : label is "42075171A10554600B3E05266170C1C08D13D1853DD28890B98AC2BD0712800E";
    attribute INIT_2A of inst : label is "6B30E18EDE2656199B9850E7E28E8CC4603FCD3F84FF7A1CD0A37457FB01B721";
    attribute INIT_2B of inst : label is "8465288CF738C06C5D9C4195F0D3DC081DA476374B0D84760A2D1372488980F3";
    attribute INIT_2C of inst : label is "20840819A28140BDF20C9081A4808E811C20C47402AC2293C2C702DB8C8CF06D";
    attribute INIT_2D of inst : label is "224A90D13468C71356B074536024831930904C71AC8C045F00142C4A102C3290";
    attribute INIT_2E of inst : label is "4514596520304B47E8E39B5D75BA28377C661CC1CFDD8CCB510D766D73319565";
    attribute INIT_2F of inst : label is "90E35D6F53EB8818186C415DCC32B34C24C1109D1C9547898D451345072FD5D9";
    attribute INIT_30 of inst : label is "96C4CDF3E4301EC4C1DE77943B76BEAA4CF40CC9954C2348C0F773499C4EFC22";
    attribute INIT_31 of inst : label is "89A4CE396465B8C0D606799AB0C24A2025C89605DEA873A955750026A26FB969";
    attribute INIT_32 of inst : label is "2B7068CC9C83610F9CE4610BC297928A3366A4AA21A877B49A91A8468B6C6C1E";
    attribute INIT_33 of inst : label is "8217A8DB25762E4018003044A95CB1769B748C6CA82A108217170F10356C664D";
    attribute INIT_34 of inst : label is "7E06DE8C3319B372641D24DDB184BC85CD68846668B933882C67492C33AA44F3";
    attribute INIT_35 of inst : label is "45BBD36BF4AC3F40ADD736D9D9C14FF4CB27143CBA5BA5943197CE319282D1D5";
    attribute INIT_36 of inst : label is "B1F24159E62EE3BBB3CCAF3C22AE3A327A647D7B819A13D3A13BF93BA75BB593";
    attribute INIT_37 of inst : label is "B371CDC58A86C8ABDDD3774D23277ECA94DD4E9675177B098CE84E846E631EBB";
    attribute INIT_38 of inst : label is "8C9DACEBE826922AF7050D8C37819763858D45ADD2F473E88B6715A30978F2E9";
    attribute INIT_39 of inst : label is "CDC526BDD7A168802A89D15771B2F3A24D14227F600030F0002AC505F5F64FC4";
    attribute INIT_3A of inst : label is "7FB87C8C0E30DFBA7DFFFFFFAAAAAA626AF7B6591F925F5FFFFFF7F75F575F5F";
    attribute INIT_3B of inst : label is "08A282BD3ACC092EFAE63BFDF43E0F868EEF6676DD2F1E9DE7B5C7E73845D459";
    attribute INIT_3C of inst : label is "AC8C0726A4D49CC10534216C8C238F48DC7761866646CF6D9E730D31CB927973";
    attribute INIT_3D of inst : label is "50111850CE48533204224805B6B49D19C4708178608AB2FAAFAFEF3FFAFA7AFA";
    attribute INIT_3E of inst : label is "8BDBFA742CCBAAF2E4DF7FD3FBA6AAAABBF5FF7F7F575FDF95ACEFFF3E158D5D";
    attribute INIT_3F of inst : label is "BAF1E7FBEA6CE3A97F3BCEF722D8BB95436B916C8FDFCBC3B7A9B85999A65B5A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "27D6DC9349446F079A39E00F0008A8FC0049D8416EDF62079451AABA5AD86CA8";
    attribute INIT_01 of inst : label is "733AD613689A9323322662305403246642BBB12B28292044D6783CF0539D0DC4";
    attribute INIT_02 of inst : label is "6204E200E73056779404252A4D5036C5188C13024526801CA0404CD820CE6486";
    attribute INIT_03 of inst : label is "C3868C931D657614338085CEF75C583338C1830988C324401100C384E33331CC";
    attribute INIT_04 of inst : label is "60B8667866559A45E3C3322E150F14253D4EF3DD6D91111710F5AE3441070645";
    attribute INIT_05 of inst : label is "0E45CEAC11B444E63F2DB32A4E6D191B73066C14E224931223A6E19E2E278B26";
    attribute INIT_06 of inst : label is "8820CAE754545C4C97FEFFE6F2B71A11020026F74A2518012B0D6DA07813C23A";
    attribute INIT_07 of inst : label is "000818A503900155000080005501540020EA38A289C7DC61A8888A229A1A1818";
    attribute INIT_08 of inst : label is "018949D020024A4360710430020A0A081E00F375A00041851842301800010300";
    attribute INIT_09 of inst : label is "8C8A68CB194A66093808D10C4C633A56501100DA28474CC7324CB0C2072909BD";
    attribute INIT_0A of inst : label is "0800228850404111022800024105500F8DC2B708582340ADC262A06212230802";
    attribute INIT_0B of inst : label is "CCA0DA2248812489E9BA6E93CD72539292AC800222A0A000A0080000228880A8";
    attribute INIT_0C of inst : label is "509A5A79149B0F1CBA90BC264D3617336AF5D2BCEC4523C4FCB87F53D645B9C8";
    attribute INIT_0D of inst : label is "19306251196905869C2E6C550A7A717A7411B288613811123D70C5B90809080B";
    attribute INIT_0E of inst : label is "5A20C608C025656DFA8F1676454657562CC63A9621266F0C9466392C14B2B0E8";
    attribute INIT_0F of inst : label is "898B03631594544633F14C60965010C2A20C631AA4E6A808E1893183208AC0B0";
    attribute INIT_10 of inst : label is "5B56C1CA1218B599B95494944586160E3831D09F18038B271831D1CC340E0248";
    attribute INIT_11 of inst : label is "FA8648C5737048612471B23B755EC3244E1103552C22704457EEF2C12B1E2F02";
    attribute INIT_12 of inst : label is "22CC4DA372D404F716A7284C5148C4CF2C42222222228BA39BBF185B80EE63A7";
    attribute INIT_13 of inst : label is "00028208641D35CD862181EB5F7DC184D3EE428040A80A628800A20A6C880B2A";
    attribute INIT_14 of inst : label is "2EB1283103443969D9AC1BC20E2A181223762231F908F90868386839F2FDF0F5";
    attribute INIT_15 of inst : label is "48514051D90650115A0462409826DF12DC4C5AE0A71F6DC5CB18AF1804973491";
    attribute INIT_16 of inst : label is "12312007D3B54819804A9A81431650508998A622A00808A082EEE08309E6F275";
    attribute INIT_17 of inst : label is "553A808051B400852A08DA2A975D65E51C2002096EF343E4FA10F7BEBEB23131";
    attribute INIT_18 of inst : label is "9D468C1310A16A57EA5E8CAF4A57855700105010242DA38F30D967C62E41D509";
    attribute INIT_19 of inst : label is "51DC10F4081A79C67353CC319A68A1870DC630B7FC824AA35C5046C4137CC5F6";
    attribute INIT_1A of inst : label is "4C3536299CE18941122F286A13AF7336BC03B440B844B043BB00B43604C0B138";
    attribute INIT_1B of inst : label is "A3845162592572FAFC064B16D6DD65DB84E298F2C922A2A613ABA0E386D8B1C3";
    attribute INIT_1C of inst : label is "8A16A280C00540104BA8A04A255C5F2A72F078F02DAC31146AD2309035393F94";
    attribute INIT_1D of inst : label is "12DA00120082C442801A081A030301A00052E2840200080000088020820A281A";
    attribute INIT_1E of inst : label is "8B880430555511458E38BC04110C1022208E80A9000240A00020040A0A868080";
    attribute INIT_1F of inst : label is "83CC0811002000201A69A3E201647C4628246200A40288200A8B00442A313926";
    attribute INIT_20 of inst : label is "4E71C0D442C6F59ED2D14C688B8D671C9BDEDA00D94D11225ECF88F24804938C";
    attribute INIT_21 of inst : label is "C8B04EE4D77D3F5C0973D24473737E185C5DE4A7A46D84670183063E1B0AABC4";
    attribute INIT_22 of inst : label is "931803C1E237EA050B4CFD4A58541014CBFC201BABF9458283082222CB319008";
    attribute INIT_23 of inst : label is "1681E20A078524974421A136169995C125A761B12CEEB0D1089C2CB04636A102";
    attribute INIT_24 of inst : label is "EAA7689F5E3C5749A8D78D28361D2E453605964A831D734BCE30F315976D9C44";
    attribute INIT_25 of inst : label is "401012880580A30170B1CD3C1255D8BB18F110962E4FA38D10D91A5AA6AFA90E";
    attribute INIT_26 of inst : label is "231CC7350131D0657338C1D5055100018280000280000000820800220002000A";
    attribute INIT_27 of inst : label is "9B2EF94A4C244824B1AC10054000D45DABB22EC9300A028A664302AE42FA6C36";
    attribute INIT_28 of inst : label is "6E061B40262206215140CB32C80A0A0C5166416E8060449F66CB4AC82D684645";
    attribute INIT_29 of inst : label is "BC4207FA9AAC8C208414016CD88EB76834124501A4710602F4261B30148902C4";
    attribute INIT_2A of inst : label is "6962E18F8441B4506A98EC53659244B88B710F63252CA3B1A1C6E05035410E8A";
    attribute INIT_2B of inst : label is "08262CCA179403209C48018B69E56C93044811A7A26C68AC1C0D1688FEF8C0B5";
    attribute INIT_2C of inst : label is "54639ACC9C31EB2E8E5CD1DD6402421CC861CB1B8534076DCD4E31505C544315";
    attribute INIT_2D of inst : label is "563E6AC6E84E7309633A13DEC8465BCBEDF63A328685152741C1383981155764";
    attribute INIT_2E of inst : label is "E38C38C3733232331916694D88C5458410CE1CC12E223F8BF2AD080331222C43";
    attribute INIT_2F of inst : label is "00F3E20C2599CCC188E2A2DA670635D7E33809CA6807800A8A4C0E0696738390";
    attribute INIT_30 of inst : label is "C788DA36D2074E0BB9B0562C0962D674847033C023944793D9E12B5B8F884B8F";
    attribute INIT_31 of inst : label is "B3C1D9152A227988CC3810049466D40344C5AE43132D6D4BAFB7936E16652045";
    attribute INIT_32 of inst : label is "3B0819931635B830816312C6952ACA9CCE4083522E44A8C1022E6C398AB33320";
    attribute INIT_33 of inst : label is "0CE1270259DB9466C2BAD818507F5E0F0423331539B214C4C0405AC5C2933130";
    attribute INIT_34 of inst : label is "700858D6B99B82120562C85334496942C284C2372E5B8D8BF6480AF48D80956D";
    attribute INIT_35 of inst : label is "88B7E6ABC012175C4822C24B094730414CC2EA0C5C9B499B902C36494F848E10";
    attribute INIT_36 of inst : label is "91D99A66933CDB76718C7F18F38DD7233A19A7310998B955819D499D5F115D9F";
    attribute INIT_37 of inst : label is "E447111C6669AEEA91144471BABAECEC85467F5659D191F52E60660642E709D9";
    attribute INIT_38 of inst : label is "1C51A13DCEA3E941F47171142B3CAEEAE91161FCE4F9E7744E046195FCB1E674";
    attribute INIT_39 of inst : label is "5051209C04825249503053540A04D95E50F3569A15450505504290500F34B1F8";
    attribute INIT_3A of inst : label is "024BA21AD92E1444A800000004040068010330414082E0800000000000080000";
    attribute INIT_3B of inst : label is "DA02624E516552B100709D4656551547277188988426B0EC8C34240EB873E7B4";
    attribute INIT_3C of inst : label is "00000259032A2E0AC01130796F535797A3768DB8138B0E0AEA8C38D234428391";
    attribute INIT_3D of inst : label is "18309A18125A0C1E4800B20046457C864E10E9530D150C000000009000000000";
    attribute INIT_3E of inst : label is "56A001CA9405514428200000400C01112A5D5ED55F5D55D5400A5002B02C0A6A";
    attribute INIT_3F of inst : label is "008882020001040020AC2108C852111F4C2C3708CC09147C20056AFECB780080";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "E2B3A1F46D31E28A017DC82ACD880A50294DBDC6960B9177D356AFD10E0CDD58";
    attribute INIT_01 of inst : label is "1CFFD8B48569261DFEAA7FB3D2F1B19B6DB4751ED0D48214CCB3B75F384362AE";
    attribute INIT_02 of inst : label is "503B0DDF58A95994E15488D5ED5FCD636330EC3598F4ADE3454899A9CD391B33";
    attribute INIT_03 of inst : label is "8C3939447594CDEF44334058596767D8E30E3E3E5BACB021E6BB8C3BACA6C6BB";
    attribute INIT_04 of inst : label is "CD15011DCC1F3688767C60D0A2EE80C5201B4CA8D6C5E5E7239F48992BEBFD16";
    attribute INIT_05 of inst : label is "5DC8EB69A915EA6E0068A069EA05F58E404219839B9C47C77E13CCECDCD3759C";
    attribute INIT_06 of inst : label is "1A01031A7D7D757E00012013195992AF795113A257F15DC5751830E76E64966E";
    attribute INIT_07 of inst : label is "580541D0FB2E517650031D615DAB5D1277A0611D9190A126D140CD03AFADADAF";
    attribute INIT_08 of inst : label is "54F4FF01C0AA8A835045F5CFAB2A67A415E34C6447B117B0AD51D0D98DFD3700";
    attribute INIT_09 of inst : label is "2999C41E8138CEE313138C118F8E8AE8348C9553D1B17A3557396F4DC7F5FC10";
    attribute INIT_0A of inst : label is "1A00C20843484811A0000030C058D015F42F51BF42D529546439F4B9466575F6";
    attribute INIT_0B of inst : label is "33074DDDF312CF331445114C378CEFEC4D7128330C004000684A300343829040";
    attribute INIT_0C of inst : label is "5779575486AAB7BC557C0832B4FE80884540A60A1D18C72FE0769AAE253A4633";
    attribute INIT_0D of inst : label is "C4B5F5818887670EF1D91B5CABC5C7D52B66FDD9C344C46B3875C09474B075F5";
    attribute INIT_0E of inst : label is "340FB68046578FC78F1353039E78F8F919B6E9C3653B19397138601970CEC719";
    attribute INIT_0F of inst : label is "F6C6442CE63FE7F9E42438ADD8FD7C7740FB6E4E6719232D94BC62B6E7DCAD65";
    attribute INIT_10 of inst : label is "567BD4D976780EFCBC79D1D9281DBEBAB3FDF78B43EE7FDD03FDF6BB9EFF6B13";
    attribute INIT_11 of inst : label is "D150C9A4CACC3CC7A8FFF4DDD87A32D2D9D9AE50D7C8312E82C3EFC68FCDF33C";
    attribute INIT_12 of inst : label is "119810BE915E4E59625077BBFFF73F75188FFFFF5F5E469E2C424936DF392EFE";
    attribute INIT_13 of inst : label is "343F7DFFD2679A6376FD3C1E259E27710491677F6FD795B7C655F195B9DE76FF";
    attribute INIT_14 of inst : label is "ABB439BD688294D49450160167BE4E0EBB1EBA0DF5F0F4F0E5555545B3BDB3BC";
    attribute INIT_15 of inst : label is "C57CE5F661BFAEE16FD487CD39C6725128C85FD41925C294EE5DB811F43B6DC5";
    attribute INIT_16 of inst : label is "01E671980F0FBF6D951D46D47DBC9E9F9E2B631F1CD1C747919B8B911EF3A580";
    attribute INIT_17 of inst : label is "824FCD776F0F77F6D1BF8B664924924204DC6E7FD1A494A7AE7B00E94941E6E4";
    attribute INIT_18 of inst : label is "4039405EE677DB5E4DC01D582AAE0A4ECAC9F9DA9BD8117D53864040997422F4";
    attribute INIT_19 of inst : label is "CE30F30BE671C71C8C1638F2299347223838C3620817035D315D2550B2D37405";
    attribute INIT_1A of inst : label is "10C24B462641758FF6320704151591D9E6DCED8CE598C39CE92E40C1910F08C3";
    attribute INIT_1B of inst : label is "DEF370B5631F91548099B6281DE19737390D679F2E2483F0E4B4B30CDB8DE00E";
    attribute INIT_1C of inst : label is "5D5157557BEBAEBA1455D5158AFAE8DF5D57F757F77FCDE69F89EF524167E271";
    attribute INIT_1D of inst : label is "55C57747AD7D7EA85D475D57FCFDEB6B55DF5D51FFF5A7F5D5F77D5777FDD5E5";
    attribute INIT_1E of inst : label is "5E3D5345EBAEBAEB51456DD1BAA2AFE03551D5D4755715A7D755515F55D1D561";
    attribute INIT_1F of inst : label is "56B2C104AACA2AC2451457F7AB8AFEEC7578175550175D755B7C5559FD646451";
    attribute INIT_20 of inst : label is "98B3ABC1B206FD3647DA29D37B6BCF6A9E19BC27A07FED931BDCDFE134BC6767";
    attribute INIT_21 of inst : label is "89FD51503B83C8FEF8EE6E7EB5CFCE38098847173425F42307CE38B399B3642C";
    attribute INIT_22 of inst : label is "C875E616591011FD4400A8B5A7FFFEA152ABE446B18E0211063777771CE4E2DD";
    attribute INIT_23 of inst : label is "C3B4A7B3985BDF381234E4E29EE6421E78F11CE4B31B4F04C16BF9E16940BCCC";
    attribute INIT_24 of inst : label is "A3A82D60AA4E27332F02C87B88BFA2D96114C3CE77CD873F93556418619E69A4";
    attribute INIT_25 of inst : label is "C0900D15C2C2634775B49B1192CA7A912C045C939535473DC33EDB5D16554CF7";
    attribute INIT_26 of inst : label is "DE0180612EEA2C9F84630911355D5B4732155540B555555060040100E8B2E0E1";
    attribute INIT_27 of inst : label is "4E5B8C176EB5E4D4E4989A78B77F7EA76467F594F11F47D9BB24F5D96DAF9140";
    attribute INIT_28 of inst : label is "61015C07BE033E89293DDEB5D94141CC0D26CE7839C3046F4BDE07C9FCBB0515";
    attribute INIT_29 of inst : label is "B0C8CAC7380F2EAA50F096682D2E8ED97D7328963285D7E644E95EC1C03BE691";
    attribute INIT_2A of inst : label is "042DB41B4DDF29E224E591969E596F16962E583EF072C7CCE4C311ACE00E519E";
    attribute INIT_2B of inst : label is "5910530778776D96ED599836810686135119445B95B979F8D4F363D72D010D60";
    attribute INIT_2C of inst : label is "19D65DEDAAD26E02E01DC6C0C71680A8C97836EE66E3761E3A30EF3D2323AEB3";
    attribute INIT_2D of inst : label is "1289E398293291AB948EAE381967A96100E28F437978C352CCEC5775196CA197";
    attribute INIT_2E of inst : label is "8E38E38C9199919C54D32618336EA38E61104D96F1B66F1006D351964045B82E";
    attribute INIT_2F of inst : label is "2786BE47CF5262779F1B378F9884C618AE6A6CDF7970BE56DFB0709AD324D4C3";
    attribute INIT_30 of inst : label is "E3DB5E827EE7AF379CA98329C3C5CDCA5179F6EFC04A2C43BCD63E56BA6287D3";
    attribute INIT_31 of inst : label is "36C8DF8E8A8AC51928B18A3636EA3C47C9D07CCE295D9E35FADAB65AE5208215";
    attribute INIT_32 of inst : label is "C559CAE6A9D257CF866C0F81D3D3E576B0940C2079B8D72E505918C640C6C6BC";
    attribute INIT_33 of inst : label is "B9AD501116674E91B7E79A6349D565F542FE6600CC49F10395B5A5BA35E6C0C7";
    attribute INIT_34 of inst : label is "71791FD1926370C41B6D09368EB5C16A56C1CD30D48E3572F2C4A7E23574769D";
    attribute INIT_35 of inst : label is "8715A583E8A6F7F00567571E2B3E8CA30DD7E5FB8C413D7FD228034639747FF6";
    attribute INIT_36 of inst : label is "115DD377C77EAAAF51045510F7EA877792DD579181B831F50115C115FF31FDB7";
    attribute INIT_37 of inst : label is "37745DD1AAB7FFDD5DD17745FFFFFABEB7F775F6FDFDB1DF04704604E0E58579";
    attribute INIT_38 of inst : label is "DFDDBD85F6C4A0E8374505DDAAA0A0A3C5DD0D6BF7FD11F01B775D058DFD10F1";
    attribute INIT_39 of inst : label is "B7B773A58EB9BBEBE4613402B9667BFDB7EE12B97DB5F5F555555555F5F3F7FD";
    attribute INIT_3A of inst : label is "F13D934F75D4ACEE95555555AEAAAB823647671E1185F555555D555555555555";
    attribute INIT_3B of inst : label is "4F3440336ACBFF1C65316819CBECFB3D5A1670671952C3B9B34D4152CD94B9E5";
    attribute INIT_3C of inst : label is "5E3E2726EDCAC6EB856761358D6BD013F663D8BDE37DF4F3FFC8B3CE49BC7560";
    attribute INIT_3D of inst : label is "ACF1DEACC4F2FDBC7C6E9F15C9E9C02F33FE5E4675E9BDF555555545F5F5F5F5";
    attribute INIT_3E of inst : label is "A76564AF9BA8000C11A0028400515EFF55D57B00A0555D5D55D625507771F63E";
    attribute INIT_3F of inst : label is "558C720600C22C0320C3E4EE2799DDD4195240F1D1165904F65A7337B749C545";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "0809027E3C2F90D521CF35E13931530B27E32BBC9204980452FD050010128150";
    attribute INIT_01 of inst : label is "7C996B9C9C6DA640182A841B17F0B756EF5A8300B8990A06771C9D75B36CC822";
    attribute INIT_02 of inst : label is "ED489112AD22B40C880D53100BB054B324492240620DD03440D5089CB08BE6CE";
    attribute INIT_03 of inst : label is "12484975D10CD11B005C30C844D0D2EB0092424BAC826003424012488262255A";
    attribute INIT_04 of inst : label is "0EA68C2ABAD84484B83CC2CBBEE848B08AE0EAB99CC96BA80B7FA2BF39999F0E";
    attribute INIT_05 of inst : label is "71973E223441A59B2A820281A4D0E41566F8A37D28B0EC58CDFD1327B1C8CF20";
    attribute INIT_06 of inst : label is "00807100606068691001A00A04C84B107D4136B76A0F9805783D69AE584D6A5A";
    attribute INIT_07 of inst : label is "F087D01592C20063D8211EC118E30802A8A8073039686880A060C1832A0A0A08";
    attribute INIT_08 of inst : label is "A4B02AD805EA808080908210082828AB6AB0426253C00891ED91400381D03C0C";
    attribute INIT_09 of inst : label is "688E1B4F693644D9434356423D642153C431242368806C948D5E70240F2C2B2D";
    attribute INIT_0A of inst : label is "7FCCFE9FBA8C9D28F2DB6EBEA1CB8BC61FF4FED31B665DBFF793DF938C5F7FDC";
    attribute INIT_0B of inst : label is "ABE3E7FF002020C2F9BE6E9B4A30AA6398FFBCFFDEF3DDFFFF5F3B6BFF5A3AFF";
    attribute INIT_0C of inst : label is "062906059CC094B2005044E71C560AB6117656856DACAFD5E4796842D5A5A101";
    attribute INIT_0D of inst : label is "32EF04CA6E28A70681ACCC4DC12A5D4AD150F4EB0A408360210091C521C53000";
    attribute INIT_0E of inst : label is "186E1689209D4220BD0BDC28D34520242216A22963A6D313C8454D3369384641";
    attribute INIT_0F of inst : label is "6808EAC48003E3F5AAE2A2BAD028DFE286E168349A021B422EE0CAE809E03AAE";
    attribute INIT_10 of inst : label is "68C07260A98A518B56C7E3224D574BF53BD5E4B908CB255ADAD5E4F25ED3D899";
    attribute INIT_11 of inst : label is "BAFA3667938C73901317263B9C5413CF233F2450B1A53C195C107CAC55038AAF";
    attribute INIT_12 of inst : label is "88099190638C0846E7156108CCBE8FEAC192222AA2AA107A68555D6630998A1F";
    attribute INIT_13 of inst : label is "4140430CBC9D8DE15D93725B5C71C8AE055166665CE695A6A4D1A8353068549A";
    attribute INIT_14 of inst : label is "1158808B55D7189B3A031C830ABBFBFBEA1EEBAF190319B040545154024C024F";
    attribute INIT_15 of inst : label is "6FD64F5C3677FE64F6D6CF8D459B21DEC333643C2E2B8B07E4920288E85C2AC9";
    attribute INIT_16 of inst : label is "214041B14A53C119C15806456ACDDA5AB749528A020A868AACB552ACAE202075";
    attribute INIT_17 of inst : label is "D7085908D99C10BD5366C965F6DB6DB67054EA8A2820F1C002A41430B0A1E0A7";
    attribute INIT_18 of inst : label is "02E50099477C405900401C102008100810514115466DAC2B96C615370B01D701";
    attribute INIT_19 of inst : label is "D24DB4CA889A69A78BF269B7D84A221C0049B4B6A412C7D30408DE0CD5145DE0";
    attribute INIT_1A of inst : label is "12B2FEEA641740DACDCFAFAC67938055AEFB4B3BCBD3CAD84FAECFCB110B8868";
    attribute INIT_1B of inst : label is "5C6B89EF5212C9F00384289717B305D6F32FBE38A8F31267CA2A1EBCC18B681C";
    attribute INIT_1C of inst : label is "08040202D04450004100804020100A807870D2D20504038046D9B4426F2EA852";
    attribute INIT_1D of inst : label is "1090201202F04402081208130101000100820814020548208888800082082010";
    attribute INIT_1E of inst : label is "FAB77BAFEBAEBAEBFBEFEB6BB2A2B90ADBFB3E1F7D1D3FAFF87F6BEB7FDACE9F";
    attribute INIT_1F of inst : label is "98E2D888AA82290AFEFBFEBDAB8ADFE8DF83BDFF8315577FFEF6FBF36B6E2E1B";
    attribute INIT_20 of inst : label is "E31CCF62D44BA263F86AF36E700C1BF3FCA2CC0E5907EB906570324E1A126D8B";
    attribute INIT_21 of inst : label is "411AE8CA174CDB8F663AF132720F9371A26525ADAEE2EEE8AD68E38992B867A8";
    attribute INIT_22 of inst : label is "54013880ACA54722B3BCA8C4080002C0A2AAB0166CEA34933640ABBA85D554CE";
    attribute INIT_23 of inst : label is "46B5EFB3ACC0D0698A35ADE64991F34979B053A478A9A2852354E9AD52A1B464";
    attribute INIT_24 of inst : label is "1817CCCC5437B8A6C799A0C3FDA7319CCC26182068874C7431CE0E782ADB239A";
    attribute INIT_25 of inst : label is "BEADBDA376F717548D5821A75E9903E68CAF9EF91F2F0CFFDAEFB5F6ADAA0E4D";
    attribute INIT_26 of inst : label is "742709E5357350B42000919921041C02001FFFC01F5F5F5040040000E0306001";
    attribute INIT_27 of inst : label is "6AD2B662EBBCE64CA6613441C100DD577AA0A0825B7FEE2BE745DCC8501B2304";
    attribute INIT_28 of inst : label is "21C1CC74965B76CD434EEA2FA01A9A75532D26C5332A8F4BCAE472EBECA68C9F";
    attribute INIT_29 of inst : label is "D12743F4197D82704925600D478877143E1141E014131F621C218E58C74862A7";
    attribute INIT_2A of inst : label is "3BC58AE82DD4451101AE222A0028AC0408C6E6D88AE17C434E398985681AF86C";
    attribute INIT_2B of inst : label is "922AAA9CB4303043267322F4C1AECE12B2228C691A0B82B38EB08900837358EC";
    attribute INIT_2C of inst : label is "61B05D980440251199292499E580CA30991C73ABB176338C4945BB6494945BB6";
    attribute INIT_2D of inst : label is "32719183502EC23976165249242DF35B89AAE3A35554644D26BD87A6106822DB";
    attribute INIT_2E of inst : label is "34D34C32080801857F9D03BA337E328AAE22C68AC2949406A8B0D1082C62E238";
    attribute INIT_2F of inst : label is "85E8114C91130013FF22AD25CCE04D3C308C4735513D1AC4A4B67B14192E9A4D";
    attribute INIT_30 of inst : label is "3863F4682CE13F74220B9812EE46CF0163F9DCCDC72DB761C73A87E8B84DA69E";
    attribute INIT_31 of inst : label is "9C2E604192939C71E3939AA6411F4745AA3A8E8A265296AF00380EA2CA2FCB87";
    attribute INIT_32 of inst : label is "812B566357BD8AB2CB5C7689F38EB288A043520D39558A920D19553BD5822663";
    attribute INIT_33 of inst : label is "6CDB562CCB1A737DEDB6D6E4C20ED2AAD912226169E825A580E0F0EFC0033731";
    attribute INIT_34 of inst : label is "CB82F121C91C3DF19CB780AC53F21453FCEA0E8E62831A78436AED431A785F86";
    attribute INIT_35 of inst : label is "EBBEFEEBEEFDB7C6B74938E1746165D4E37C37E28045A3113B12CDB036FA33BC";
    attribute INIT_36 of inst : label is "560AAEAAAAA04710157501572A447AAAD7AA0755CD5655516D513D5121552150";
    attribute INIT_37 of inst : label is "8AAB2AA21114AAA82AA0AA82ABAAAC54480A840552A2D500B55B55B57F59DA95";
    attribute INIT_38 of inst : label is "AC3AA2C57974A1D5CAA92AAE2062A1E072AABA1CAABA015118AA914502AA6150";
    attribute INIT_39 of inst : label is "444D85A60FC0B843A06B769CB600F15A44D236C93DB0000000000000002EAABB";
    attribute INIT_3A of inst : label is "57BB79A49451CEFE7BFBFFFFAAAAAA12A4E42AB88B869F5FFFFFFFDF5F5F7F5F";
    attribute INIT_3B of inst : label is "E1E055E16A7BFB066B1B20C3ECAEABA4C830ED0E43910BC231C349B1073E516D";
    attribute INIT_3C of inst : label is "0404981F02E97820D8163364CD33CA8CAA62A8E552730C20504B34D2C8438081";
    attribute INIT_3D of inst : label is "58705A580A58229E184ECF605251486743AF5EB410680A000000001000000000";
    attribute INIT_3E of inst : label is "945FFF747D8BAB18BFF8BEBD14AAAADFEE042BEE4ED6DF4FDFB80EF2364BB810";
    attribute INIT_3F of inst : label is "FF3FCF7CEACAB3ABF73D89414DD7D78C53D7CF0FBC47931C6EE84519FD277C6E";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "6FAEAFF31D17FCE539EBF86F5DDDF3E9D0FACC37239C6A4C54FF003F5A9B41A0";
    attribute INIT_01 of inst : label is "F7D8B72F79F697F4A9AFE8983D54755FC62ACA836A7BACD8F739A874C7991C43";
    attribute INIT_02 of inst : label is "ECDEE22227B73B663EDE24C6F9120853798F3F8E6F7E831B0DE27EC6334C3EFD";
    attribute INIT_03 of inst : label is "E7DEDE8A5964EB297396D2DEB7E8C955F8E38FCBA3C3BF537798E3CFE7BB5A4F";
    attribute INIT_04 of inst : label is "99A2FECA179FDC4F3B3BBCE65578095CE27F25867A1B8FAEC988162C52120718";
    attribute INIT_05 of inst : label is "6C92B2BF57D559F3C7EFADE8F1B555678DDABE65FA19BA26AF3E96AC81DEAF29";
    attribute INIT_06 of inst : label is "EFFE325B8B8B8B9D9D54554C3F23C3A2C3AB0F8E7E4BDB014F82A6E3FA0AE8A8";
    attribute INIT_07 of inst : label is "AEEA9EEA4BF8739CABBEEABEE700F318D5CBBF0825BFEFD73EBABAEED7575757";
    attribute INIT_08 of inst : label is "A94BB6EFF55D7775EEFBAABA971DD35BF858E3BB94C14F90E2EEBFEE5A0E5ACA";
    attribute INIT_09 of inst : label is "AFABE36EE9D577558F8FCD8C766F3577ED38889D8942FAE6667DDFAABB37C7AE";
    attribute INIT_0A of inst : label is "AFBFBBBE20830204AFAFABAB1AA22C8C1FB46ED15FFE4DDFB747F6C75B2E5C57";
    attribute INIT_0B of inst : label is "BE426AEA08A42B8ACDB36CDB8AE286EEDA3AEBEE4B0F1B4FBEAFEFBA8A1F0A1E";
    attribute INIT_0C of inst : label is "9BA69BBA875B724BABA9AC3A516F3746793F982FDDDFD727C97B43CF05684F8A";
    attribute INIT_0D of inst : label is "735669F8EEFBBBEFFE0ECE8AD1B96EF3B3623D3269EE7F7FB67C66EACE0FCA8A";
    attribute INIT_0E of inst : label is "1566EE778BA96200F54F7F2A41062626DCFE26AAA90CBFCF6EC079CE6EB0D8E1";
    attribute INIT_0F of inst : label is "2A37A3A1FD8BFF46FABAEE76820ED358566EE3AC9645F8C1E9CBB9C706A5D6FD";
    attribute INIT_10 of inst : label is "FBCDEBF0CD377D373ACF4E8E99C6C53598ABCCB03E23E23AC9ABCDCE6D1132CA";
    attribute INIT_11 of inst : label is "F7723EA8F679BD7DDE29A62D781986D5BEB6551511640E61BB17B2A3629B8FCB";
    attribute INIT_12 of inst : label is "DCC6EEB17A4DC4B7DEAABA3A04010053D676AAE8AEA8B5AD93AB6F6B264EE7AA";
    attribute INIT_13 of inst : label is "9B924B2C47FC238CCE338CA3F966F69CDAEE9F9862288A4FF2ABBCAAEEDE0B3B";
    attribute INIT_14 of inst : label is "CE2F0201059D78F9BAAC338C37FB5F5DA842AA08030C030EAABABAB805010501";
    attribute INIT_15 of inst : label is "6FD74F5D11D4776EC6AE12335675FD8ECF6FFB378278B859C3AAA72013E0DC9A";
    attribute INIT_16 of inst : label is "F6B3A33213616BA9AAABD82A516716D42A90B6CD6BB4B2D20DE2A30D97B7422A";
    attribute INIT_17 of inst : label is "28BEE3BF78A6BBFC50C8F8A3B3CF3CC1F828C833B744153970392EBDBCB6035F";
    attribute INIT_18 of inst : label is "4546EFE393B9FDDE6AC1ADBDFC5EFD57FAEBABAA38BEAC013CFBAAF6F2FB5D4B";
    attribute INIT_19 of inst : label is "E78E3CF493BC71E62353CE39BE32E2F9898E3D3FFCFE7CF3CCFB586F075F40F5";
    attribute INIT_1A of inst : label is "5E76763A9AED82E8AFFE1F1DE7E22655B62639F63A4F19127D9D963F45C47B79";
    attribute INIT_1B of inst : label is "33AE9F6678E067BEFF577796823AE0588FE2CCE6D746C21A3E7639E35F793BD7";
    attribute INIT_1C of inst : label is "A7ABADA655D5D5D5EEAB2BEE55654957FD57F05ACD565B267C673CD975DDDFE5";
    attribute INIT_1D of inst : label is "BE3F8EBCF7D551D7A7BCA6B4D5D5D5D4AE2CA6BFE8FBFA1AABABABAB78E2CA6A";
    attribute INIT_1E of inst : label is "EB2B3FBFCB26BA49BEFEAFBFB08A8A02EBBF2EAB7E5C7E5AAAAFAFFF6B9FCE0B";
    attribute INIT_1F of inst : label is "A32E70FF08A88A80EFBEFAD8218A020C9FFEB9BB7E58163FEF62EBFB193D4F1F";
    attribute INIT_20 of inst : label is "0F3DC8FE498B51A4DBB9CCBDE5D8E5A37BCEC0C9635B1F38F8ACAE946B339A13";
    attribute INIT_21 of inst : label is "222AFAFADF505CB5DF88C83C64FF74D6EF6F125A092229AB2847CE6C5ACEA6C3";
    attribute INIT_22 of inst : label is "1D7A6FEBA6BDE47A335DBEA54AABFF6DEFFFCBBBAEF745008B8A8C8DEA8A08A3";
    attribute INIT_23 of inst : label is "7E8A82083E893CDBEF0AA2BB368AD307B7EF62337F6E3A5D70AA8E7DC79A9502";
    attribute INIT_24 of inst : label is "BFBAA8ABA9129D95FA3EBDA8D463490EBA9FBB2AAC1E7F0EDE6DB797B672BD63";
    attribute INIT_25 of inst : label is "AFAABBAC4543E719A72FCF090F0F467522E60C7F0E55EA4F38C52CE92F55E4AB";
    attribute INIT_26 of inst : label is "6FBFEE8942E1146CF379E6ED0E11A184EFEAAAAF8A0A0A0BAFABFEEA1B0E0A3A";
    attribute INIT_27 of inst : label is "6799E6B55D65D0343FA678CD2BA3C57993F98DE9B85F40E03C3AD28FC37AEED7";
    attribute INIT_28 of inst : label is "3ED68FF64FF46FFECFDB27DACCF6F671F7EE6786B6A95FE399E6F5F22FC95F5E";
    attribute INIT_29 of inst : label is "66669FE29DAAD9452F0A0E4288D3C62C70A1D90EBD7F1F23FDBECDF85FCF23CE";
    attribute INIT_2A of inst : label is "D1A177DFE550F514C21CEC65A0821C0D08FDC3AFDFFF6F7ABBDA637B35D3E64E";
    attribute INIT_2B of inst : label is "26D7AAA0B43882A89CEEEDC3600CE11EAEE6BBC74A5EC63F76375FB1DE39D6FF";
    attribute INIT_2C of inst : label is "3D71FE582CF1EF1AFE1DF196171337BB7D5D87E7B78DCF6FCECB3AC8CCCC930C";
    attribute INIT_2D of inst : label is "FA0E5896FCDCB77FF5B8639FEC1E1F579EF864A02F2F3DEB625A92D3B17C5136";
    attribute INIT_2E of inst : label is "F3DF3DF5AEF00F071BFEC18DB1C4045459DE5DF396DD09AD581732AF3F2A4FD3";
    attribute INIT_2F of inst : label is "8DAB68361B89B812D9E088FFE653A9B6F7BCC3EBCA121709AEE8DE309B7FCFFD";
    attribute INIT_30 of inst : label is "9FC8FE6AF5905E6C83BB3B8FBDBE0E756EF33BC9AFBCD7B3C3F5AEFBE0936698";
    attribute INIT_31 of inst : label is "2BB7BBAB7C74F9E6CF2378CED57FD51936FBEE377CFBFA6FAFB5CAFD8FC56CDA";
    attribute INIT_32 of inst : label is "5B72A99BF60688179F63F8FE97C3DEBBFE77236C2EAABBD3DCAE2A3BB2FF1B3F";
    attribute INIT_33 of inst : label is "8CF7AB0D69BDF277FE78D8DCD526CA01BF23BFF7333E7EFECE0E1B44DF5B5F96";
    attribute INIT_34 of inst : label is "F6E67BBEDD6F9D6CAF1BA2ABBA46F014E07AB3A2B39BAAFCBF6E79BFAAF61D6F";
    attribute INIT_35 of inst : label is "37D90CB1227D9FD6AECB3B6DDDD134D56FAA962E9A5F4BD2F98DD6354CA391B4";
    attribute INIT_36 of inst : label is "2609DB77402CE9BF32488720820EB831A79DEBF21B0052021B260F26E132F785";
    attribute INIT_37 of inst : label is "4115C4451992626444551144898F84FA0157180C01F5D2C06C83C86C034218C3";
    attribute INIT_38 of inst : label is "02846D663CAB33CA250E41034D133030050544457060F8B99041566641C15999";
    attribute INIT_39 of inst : label is "9C9C2EA0D7177BCDDABAF1CE7FB74D7C9DE7FA2A99F7FAFABFEFEFAF8A14E431";
    attribute INIT_3A of inst : label is "FD3BD02F8C708CC5BCAEAEAA001000FAE5EFBAEBCBAA8A5AAAAAAAAA0A1A0B08";
    attribute INIT_3B of inst : label is "FBFEEA7E264AA7EEBAF65BFE7E0781AE96FFAB7A7E0F521FA45CC69F78F59F30";
    attribute INIT_3C of inst : label is "888883BD7FB7DF5F83B662F3350D4702B9BBE7B2AF0F9EBBEA8F3DE6F6E8BB0F";
    attribute INIT_3D of inst : label is "BCA3EABC575F5D5F6CB8730EDC1377878B833F132FB79E0AAAAAAAB28A0A8A9A";
    attribute INIT_3E of inst : label is "BFA2ADBC3C822620EAEFAABA2AA80282AAF3FAAA0A030A9A0E9ADBAD2ECFBACA";
    attribute INIT_3F of inst : label is "EFEBAFAFB0609241EADB8AE20441D5C446DC3337846EBC5F4AEBFCF3B7280C0E";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "94153D48702C02F2415D3B01A0640ECEFD8132DA04139775BB53AFFA5114BC59";
    attribute INIT_01 of inst : label is "1CB77E9C9C6BE2109680600AE0C01193E79635BCA1900A0ECC92525F2926E22C";
    attribute INIT_02 of inst : label is "32232CED4F8914477620AF29411AAA47E3B2CC37BD228D64B228D111E511A1A1";
    attribute INIT_03 of inst : label is "0C31286411C5F8B6CCBB60223C52708DC22AA63593883D0BCE3B28A28C34049F";
    attribute INIT_04 of inst : label is "4A16417DC041A2C1E44F121954CBC68B4A174C22D5C7E3E1BB930A97096BB496";
    attribute INIT_05 of inst : label is "014969EDFAA08E94634503438C70A09163F18CEA8136D1CB10E140437625E134";
    attribute INIT_06 of inst : label is "FB658BAB2525253476AA2AB3F90FAB835F1D9565787DD1D6A59A414E34C4C4F4";
    attribute INIT_07 of inst : label is "5D356F79A19A51FE528D755D7FABFD1208EBEABB38C3DD0ADB0D6431B9DB999B";
    attribute INIT_08 of inst : label is "EFAC84DFC0AFCEC269740505E2B936E6CA7B7C86AC8E093F0CC7F955EDF5F5D0";
    attribute INIT_09 of inst : label is "272268E29C31B3E4A3A137A312F3553F0F823E631E8C64F994C9B86109D9B18D";
    attribute INIT_0A of inst : label is "334C7BC8D7DC7DB13669379ACFDFF959FA77F8FD8F7F0DDA3FF715D76C57321C";
    attribute INIT_0B of inst : label is "462605458CD23B8CE7BDCF7A0CE3A92E7B9B0C91F4B2E5B3CD451A797B84FBEF";
    attribute INIT_0C of inst : label is "3503353CC0EBA3B80486BAB12082549368B3FC3A56118B28F096C7E6261F5F34";
    attribute INIT_0D of inst : label is "1B1F131B131F54370B426320A49CD28D1FCB95390BDD872B4CBEDD4625C322FA";
    attribute INIT_0E of inst : label is "C0ADA0C8B4640962152880C59E7C109023A099E064257330C2D4CB30C294EC73";
    attribute INIT_0F of inst : label is "15489A0F942CD4402EAC1EEB1091B0460A9A0E04DC14AB2783B2FBAE1CC0CB62";
    attribute INIT_10 of inst : label is "57E5640BA74807681E6429E16C5F72671B387E45518F1913BA387FE89674A830";
    attribute INIT_11 of inst : label is "EECAD244938048F20A95D694002563246D7AF8FAA4E2E62CC5EFDC5E9144EF10";
    attribute INIT_12 of inst : label is "67319D3AD85C5E3DF11256846622622422ED450564648834BAEA949F701DC826";
    attribute INIT_13 of inst : label is "363C61C684528B22629C273831CD2D07AEBFA5320D331BD41CED0733DFD04F74";
    attribute INIT_14 of inst : label is "2192191C31447C8D46FC9CE3470E0AAA10011011504050411005000444B444B7";
    attribute INIT_15 of inst : label is "CD54455456937795EDE2ACE90D52A753EAA0C5FCB3694A0C7C740A995E094B47";
    attribute INIT_16 of inst : label is "6B3E6BBE8D397AE561846E7669269EDA14B92F24A4830CAD323B2D33962B1F20";
    attribute INIT_17 of inst : label is "82772FCD5A37AF47A9B313061C5147462E62F4812B0B086AA0D2C0C9A9A90E82";
    attribute INIT_18 of inst : label is "5EFF66FCD79CA022E0BAB30165A2D0FB65625361B20D16619AD542C8F8F125D9";
    attribute INIT_19 of inst : label is "5862927DE76B9C13F8FA6AB36BF47C647A609210AB3C0A596745E74BF0D86F0B";
    attribute INIT_1A of inst : label is "B0DB998711B2959BD0D52FAE9345D1A896EDCF0EE83A8B4BC42E7ACACB8F12EB";
    attribute INIT_1B of inst : label is "FE492F9D718ED958A8BF8EBA1251C4B1AA095288103AEF3EEDF5E22C3AA66A8C";
    attribute INIT_1C of inst : label is "278B8DA021A1A1B0EC270CEDC4A5D48580A0A2A82000F7BE914997125FCBCEEF";
    attribute INIT_1D of inst : label is "B5B7AF9DB70701F32E97AF89BCBDA5E127A58C0A723250F00505072578FADAAA";
    attribute INIT_1E of inst : label is "FCD7F2E269AEBA693AE2C05BBAA2A928FD7BEC147557175570F570701DD3CC15";
    attribute INIT_1F of inst : label is "CEBCC962AA02894AC5965ED7AB0AA8A8EF2119CB215E5D3E7E1FFF1D4C6C3419";
    attribute INIT_20 of inst : label is "EABA6358C6D08C22C0D36B6A912F1658ACA8FEA3782C8B800641C5F31D9E416E";
    attribute INIT_21 of inst : label is "451F6B6A26C8EAAC107EE4C54882F33EC4056DA1124D62C086FA699311A320AE";
    attribute INIT_22 of inst : label is "73DD8DC7CFB4A651CCF6BCCA6280849473FF4A0732D88B11B7B104519C4CCB05";
    attribute INIT_23 of inst : label is "A411451B122B44180BB044740C24178F184B8C4A2B11652E894971EB0FE8B84E";
    attribute INIT_24 of inst : label is "60625E1B549978EAC505D64355A9F6D149A105E46BC19463A2976863494C2A0C";
    attribute INIT_25 of inst : label is "5338513A70747E575912A29750C1388AE5FA72A5306AB4178236F3B41C0AAB40";
    attribute INIT_26 of inst : label is "4B2A9AA87BA3B48ED8C3080827DD5BE7D0D5554ED5555552DD6E9BB3EDB86BFB";
    attribute INIT_27 of inst : label is "D8FE35A56405F846C2A8C2FE7AEBE4D176A55402B937E5C3D28C79D34D74AA59";
    attribute INIT_28 of inst : label is "80A4E42DD2C57251E4E444B71D870782F800EF82198A1ED9AE57E549D4B81E0E";
    attribute INIT_29 of inst : label is "00EF6270EB5E1C708CB8A4E04E12435DBF1B72A417474C384E00E60F6261B8B3";
    attribute INIT_2A of inst : label is "4B0EBCF91D9F99A60C22172C8E34ED98B6407F54714BDDAD05200BF4EE8CE086";
    attribute INIT_2B of inst : label is "196A5190D65323D26A233F34C187C211C999263A9B7A1970808AE103A33D8B66";
    attribute INIT_2C of inst : label is "B2E811C3EB9C164E03BBE8A9CB47C4E94FEFE604D8EF28BD6878B97326272B77";
    attribute INIT_2D of inst : label is "30AB69AB7D25179C2896BEEA1D6BFA82284680499495DFC1E9EC96743B2E9B8D";
    attribute INIT_2E of inst : label is "2C32CA2C1108989266440DFA2D686309C733ABA83B2474B2AEEA81100245390E";
    attribute INIT_2F of inst : label is "2F61F4CE851A424732B39F15888687148ECAE434310EBC4645BAF2BE6125CC53";
    attribute INIT_30 of inst : label is "64F994142BC2BB731C038100C28307DE19DBB46303060E41F42C05D7F16803D3";
    attribute INIT_31 of inst : label is "9FE85985878FCD1DEABB82A043123D54EE203EEC6BDCBD01FFFFBC4FC47A8A0C";
    attribute INIT_32 of inst : label is "CF9163303C8710956628271913A14B1CD08CACD3FD12D1CC337D12C0C8E44724";
    attribute INIT_33 of inst : label is "3BA81B3253D19E86B1C70AFB5B4454214ACCC82C7CF113E1FF3F29C8905002CC";
    attribute INIT_34 of inst : label is "493914490740B8D3ECC50128D792902E64086D5CBC85335A6CE2AE6E3358263F";
    attribute INIT_35 of inst : label is "259B0CA055BEF38135BD4C277C7FC7FFA04D6E8180013F21320226CE21DE34CB";
    attribute INIT_36 of inst : label is "A0FF591D202A6D9AFACAA3AC02A6F02085349112070ADA4227A23FA21BD2470C";
    attribute INIT_37 of inst : label is "A730DCCD289E22015CCF733D888A82E0B50962EE1442920E9EBBEA9E0F421383";
    attribute INIT_38 of inst : label is "838CB1CE40A870036300488A4D353076708DA876321051989E233C2608C87099";
    attribute INIT_39 of inst : label is "BFBFA33F51F1A69852198BBB4FB6989BFEDA3487663A0A0AAA87AAAA00537A20";
    attribute INIT_3A of inst : label is "6991591541C480E8575955D5AAB8ABC07C2DA2080904354555555559555D5D57";
    attribute INIT_3B of inst : label is "8133EB9B4AEBF01A86E9EE309CC9B279FB8C2AC2902FCB351DAA182BCA8C72CF";
    attribute INIT_3C of inst : label is "2AAAAF64EC8796492D24F954E83A815605410416E5C258A0AAAAB3DC54FA7940";
    attribute INIT_3D of inst : label is "0609040640026800C204B4A5BBACC89670C2D3082C84B6F00505059730F070F0";
    attribute INIT_3E of inst : label is "05D476762CCDFBFD3BE9313CFDA0AE2AC659579313F9F595F59DC3225CDE3D64";
    attribute INIT_3F of inst : label is "553D5C34E69FEF1AC3E1541026693104FF7F5C8F4C9506A656505BF30BA55545";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "9D9CB3E86070183270CE7707E444A7A47D36BACA04D945669652AACC83CFA0A9";
    attribute INIT_01 of inst : label is "CB30C99B24D90611B08D62AF34157023A8318D3301016A06599622CADCB2B65A";
    attribute INIT_02 of inst : label is "C54C633380A3B22742C463C2C99010813C8F318BB066C36F1C662ED7F64FC3F5";
    attribute INIT_03 of inst : label is "E3CFCF5F8B244E251D4CF8C4B2CACAEA1C4343C08451204047DDC34C512B1701";
    attribute INIT_04 of inst : label is "0A8DCA2FD4D47404AD2AAA96808CD59EE9F979664E79199AA61201B6D9595E7A";
    attribute INIT_05 of inst : label is "248AA8C38F455704A8CA2ACB55515537263D085CA7800AEBB0888EC3583E5390";
    attribute INIT_06 of inst : label is "ABA2E10827252D3A9A01200B0980AA008C6A12154A0F0A1D6EB3008D40D708CA";
    attribute INIT_07 of inst : label is "A1BA9EEC82188000AC220AA000000082823F8E12314BC9009A668B9A0B090B09";
    attribute INIT_08 of inst : label is "A0AC819A15551015ACA8AEBA56ED799BE86861372C468B0DC3280BAB604A9A9A";
    attribute INIT_09 of inst : label is "800E210CA062018828089A0A73D7550F8021B5EAFEAC0613AB6F98AD09B9A219";
    attribute INIT_0A of inst : label is "42C82D858800802040BB650620820203358056011CAC42918387200728646A6A";
    attribute INIT_0B of inst : label is "AA267888845219068822A8A206418284A1349000524019120B5100501448020C";
    attribute INIT_0C of inst : label is "84838C8D00D5D195A8243013C92311A08A660C11D4ED13B0DE156A0798F12CF4";
    attribute INIT_0D of inst : label is "A28396592462B4870AE685042160E221477298190025A31B401041AF2DEB2A0A";
    attribute INIT_0E of inst : label is "75BF6FDD144E094AAA609E5E5D7A9090EF6F831F2D62AC6E3800B2EF988E8C3A";
    attribute INIT_0F of inst : label is "A0BB38C61C2C5E60A52D2BBCB0B392CF5BB6FD70CA19EE277EE8AEFD5AC99CDA";
    attribute INIT_10 of inst : label is "52AAEA23975887D8B12260E2C4FD87D21F9BA2EF2B1EC3493E9BA2A5FA0A3AE2";
    attribute INIT_11 of inst : label is "EDAFBAAC6161D3572ABCEB956060657D4AEAFE5580C2FCC8BE296EEEE3C07710";
    attribute INIT_12 of inst : label is "1058E00622C4DAB207BE0904EEAAEAA84D100005317093714AF05C186800017C";
    attribute INIT_13 of inst : label is "CB538618ACCA26AA9F6744E9892C8CAF0A08404C54641E1200FC853E03005A48";
    attribute INIT_14 of inst : label is "0E39B32D714105E78550AB2EC3E5B0E10B5E0A4F1E5B1C520FA9A500070D070E";
    attribute INIT_15 of inst : label is "C079E0F3C7B682642145A9AAD58396D525C662FA1311CE05379E2BA9EA8B17F9";
    attribute INIT_16 of inst : label is "31E670034E93204DEAC32A53620C5E581F49E280E6CD42B7047DD2054430C27F";
    attribute INIT_17 of inst : label is "7DA4D4C8F29205EE014D592FBACB2CA734709C0138D75321283DF95A9A9146C3";
    attribute INIT_18 of inst : label is "E3F848E1A129856302100822041311A18E88AC8580EC80223CF8EEA68A0BDD0B";
    attribute INIT_19 of inst : label is "C38E3CE1128820A361F38F3CDCC80849508E3C9F5582C2238B63F56CE4D15F55";
    attribute INIT_1A of inst : label is "44C78AAF1B42140072F32BAA01E5224DFC9C3E589065B71C3962E0BEC44E4DD2";
    attribute INIT_1B of inst : label is "49B268AAF0242A526DB1316898CB264B664A6E6A416ACD7FDF777AEF247A19DB";
    attribute INIT_1C of inst : label is "A2AEA8A754401544EBAA2AEAF54531AA2FA5AFAFDA786B32366019B82F6B6531";
    attribute INIT_1D of inst : label is "9A3A8AB85252D157A2B8A2AF4B4B5494AA20A2AE000AFA08A0A22A8888022A1A";
    attribute INIT_1E of inst : label is "8B0004504104104104102814102803E8648481E4104B48408F14068A00848150";
    attribute INIT_1F of inst : label is "DDABF999002003E8124923A201A02842207F4200574A0A288F8900001A150104";
    attribute INIT_20 of inst : label is "C59633E6A68119977A56276F34D673D585E72E26016431EAE8E46B7FCF8AA90A";
    attribute INIT_21 of inst : label is "AEB4C667E325095D4895AEA4E776471D79FE07A8927852FD8131A7900853E298";
    attribute INIT_22 of inst : label is "4A9D968A01900AD013B80370000007DCA80198A8698EC03B984C00105B191404";
    attribute INIT_23 of inst : label is "463CAE1B90114C188C3D8F800A0FB15D19817510604E9C702323A4B8539FA226";
    attribute INIT_24 of inst : label is "A4A2ED1A5581696F5B3E79CB37949714C7679F62D853AD2BA29B6A696B460A2A";
    attribute INIT_25 of inst : label is "220CB95600845AD768B9A9BAD10485F7E1D9DE8CB27A5C349722D394340A02D0";
    attribute INIT_26 of inst : label is "2A7A8F8D780175CCA1BCE0CD60A000082AEAAAAA0A0A0A08BCF2BE8C0B0A1302";
    attribute INIT_27 of inst : label is "892A78D0E8AC4ECCD3797C1920414C6B35F2036BCA6A0B83852B0FE45008AA44";
    attribute INIT_28 of inst : label is "034B0090E2764275818C0126E02C2C40C507002D8168CC29224AC0693478CECC";
    attribute INIT_29 of inst : label is "2327C22F89FF54608B6B4B23AF5672D43CB219CB01D34E50640B0024892340B8";
    attribute INIT_2A of inst : label is "BAC6BCF3359E9596E6AE17AA4C30452813AA68AA720B93A6273FB8A89DDA1BD8";
    attribute INIT_2B of inst : label is "4190666AD0D32B92AA6BBA6B230F23B2F66199CA97720165FDB0CC95903ADE9D";
    attribute INIT_2C of inst : label is "1CC69E880A0962310931E6008A10943D25E48B316059308D8C9B358CE8E913B8";
    attribute INIT_2D of inst : label is "360AAB0270365799B2B2270DA42C9B0A29CA08C1FEFF202E028F4CEE0118114F";
    attribute INIT_2E of inst : label is "DB6DB6D9022222A1721AE6608D68841CAB338B0C392241B8A0F08191192D765D";
    attribute INIT_2F of inst : label is "631A02BEACB28881668119F2AA4A4CB25D5627325B5F8E50631EAC887E700B4E";
    attribute INIT_30 of inst : label is "2C33B29E9D558954072ABF2E7F0105ABA44A952EEAB2DCB1277ACD52F21EA241";
    attribute INIT_31 of inst : label is "BAAC998ED2D324B5259AB6A5C7061BD4AA4C3FAB10365511FAE83749F4BEEAC7";
    attribute INIT_32 of inst : label is "0D21FCCF1A2E82AD9F76334CB18981340631635DE3D58A93CD635519969B1065";
    attribute INIT_33 of inst : label is "5DF37684C00B36ECC6D35C8CD320C8A8CD35FF320E819A0A2A4A5A45CA0F53D3";
    attribute INIT_34 of inst : label is "D931FF64F69D700341AA2B21013565726AA6A9699C5CC2E0C1A2A0C1C2EAD295";
    attribute INIT_35 of inst : label is "5561D31F8F5920330618A9EE6D79E82AE068A9AB58B10EBB962E228C69FACAE9";
    attribute INIT_36 of inst : label is "60A22088799D10452E7BA2E799D12999ED22A006FACF0E86FAEEAAEEFE06FECD";
    attribute INIT_37 of inst : label is "888AA226555C6665A23A88E2999DD53D496C9B7B22FA06F7E3AEBBEB3A3EEA4E";
    attribute INIT_38 of inst : label is "3532827645797F9B48FE5232497F7E3FD2325A7E2C3B6F1FD4C8D27E73830D1D";
    attribute INIT_39 of inst : label is "0001039CC191C180FA89949ECF460B3C81E736AF60B00A0A80282AAA0A0DAD33";
    attribute INIT_3A of inst : label is "B1D49BE3E1C6A0E99A001000000001D2904E69B4810D60000000080000080002";
    attribute INIT_3B of inst : label is "7C0A80D4C2C152202C3BE90080C8321CFA4011810043EB9B3942122ACB1A28EE";
    attribute INIT_3C of inst : label is "840410224554B2E91021516D8C6B95918876218F14F2E8D0A78F3CE42E0102CA";
    attribute INIT_3D of inst : label is "84818C84C06264B02004A4409C427D269945F4867CCE120AAAAAAA3A0A0A0A0A";
    attribute INIT_3E of inst : label is "7714838907A0AA00028987A908D7DE00B100007555005580E366000A43124716";
    attribute INIT_3F of inst : label is "459019060088088290869DAAAA6A11A402A54B18480C1C24502775244EDD0302";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
