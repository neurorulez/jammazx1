library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog_rom is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog_rom is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"00",X"E8",X"ED",X"56",X"3A",X"04",X"D0",X"A7",X"F2",X"00",X"33",X"CD",X"F4",X"05",
		X"CD",X"F2",X"06",X"CD",X"29",X"0D",X"C3",X"68",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"87",X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",
		X"EB",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"D9",X"CD",X"6D",X"05",X"21",X"4E",X"E0",
		X"34",X"7E",X"23",X"E6",X"0F",X"20",X"01",X"34",X"23",X"35",X"23",X"35",X"3A",X"04",X"D0",X"A7",
		X"FA",X"93",X"00",X"21",X"4E",X"E0",X"34",X"01",X"03",X"00",X"21",X"4E",X"E0",X"35",X"10",X"FE",
		X"0D",X"20",X"FB",X"D9",X"08",X"FB",X"FB",X"C9",X"FB",X"CD",X"8A",X"0B",X"3E",X"01",X"32",X"4D",
		X"E0",X"32",X"0F",X"E5",X"3C",X"32",X"08",X"E5",X"C3",X"B7",X"0B",X"06",X"00",X"AF",X"32",X"4D",
		X"E0",X"21",X"46",X"E0",X"70",X"FB",X"CD",X"45",X"07",X"CD",X"8A",X"0B",X"C3",X"B7",X"0B",X"06",
		X"04",X"18",X"EA",X"CD",X"CB",X"05",X"3A",X"00",X"D0",X"2F",X"32",X"53",X"E0",X"CB",X"4F",X"28",
		X"15",X"3A",X"04",X"D0",X"CB",X"67",X"20",X"0E",X"21",X"46",X"E0",X"CB",X"4E",X"20",X"07",X"3A",
		X"00",X"D0",X"E6",X"01",X"20",X"F9",X"3A",X"04",X"D0",X"CB",X"5F",X"20",X"06",X"21",X"F3",X"E0",
		X"34",X"CB",X"46",X"FD",X"E5",X"DD",X"E5",X"CD",X"0E",X"04",X"3A",X"41",X"E0",X"A7",X"20",X"05",
		X"3E",X"02",X"32",X"48",X"E0",X"21",X"46",X"E0",X"46",X"CB",X"78",X"20",X"15",X"CB",X"48",X"20",
		X"1B",X"3A",X"48",X"E0",X"A7",X"20",X"1D",X"CB",X"50",X"20",X"11",X"3A",X"47",X"E0",X"A7",X"C2",
		X"8F",X"00",X"CB",X"40",X"28",X"06",X"CD",X"7A",X"04",X"CD",X"EC",X"01",X"DD",X"E1",X"FD",X"E1",
		X"D9",X"08",X"FB",X"C9",X"36",X"02",X"31",X"00",X"E8",X"FB",X"CD",X"29",X"0D",X"CD",X"33",X"05",
		X"28",X"FB",X"CD",X"38",X"0B",X"C3",X"B7",X"0B",X"31",X"00",X"E8",X"21",X"46",X"E0",X"35",X"FB",
		X"F2",X"68",X"00",X"CD",X"96",X"0B",X"AF",X"32",X"A6",X"E1",X"21",X"15",X"E5",X"35",X"28",X"1B",
		X"CD",X"D5",X"06",X"21",X"46",X"E0",X"CB",X"66",X"CA",X"B7",X"0B",X"CD",X"03",X"06",X"3A",X"15",
		X"E5",X"A7",X"C2",X"B7",X"0B",X"CD",X"03",X"06",X"C3",X"B7",X"0B",X"3E",X"1B",X"CD",X"75",X"0D",
		X"21",X"46",X"E0",X"CB",X"66",X"28",X"1F",X"21",X"ED",X"2A",X"CD",X"4E",X"03",X"3A",X"46",X"E0",
		X"1F",X"1F",X"1F",X"E6",X"01",X"3C",X"CD",X"BD",X"03",X"CD",X"03",X"06",X"CD",X"E4",X"05",X"3A",
		X"15",X"E5",X"A7",X"C2",X"B7",X"0B",X"21",X"02",X"2B",X"CD",X"4E",X"03",X"CD",X"1C",X"06",X"28",
		X"03",X"CD",X"03",X"06",X"CD",X"E8",X"05",X"CD",X"29",X"0D",X"21",X"2A",X"2A",X"CD",X"00",X"03",
		X"3E",X"11",X"A7",X"28",X"3D",X"3D",X"27",X"32",X"54",X"E0",X"11",X"33",X"82",X"0E",X"02",X"CD",
		X"AE",X"03",X"3E",X"40",X"32",X"50",X"E0",X"3A",X"50",X"E0",X"A7",X"3A",X"54",X"E0",X"28",X"E2",
		X"3A",X"48",X"E0",X"A7",X"20",X"0B",X"21",X"57",X"2C",X"CD",X"74",X"03",X"CD",X"27",X"05",X"18",
		X"E6",X"CD",X"33",X"05",X"28",X"E1",X"CD",X"DA",X"01",X"CD",X"DA",X"01",X"CD",X"BF",X"0C",X"C3",
		X"B7",X"0B",X"F3",X"AF",X"32",X"46",X"E0",X"C3",X"68",X"00",X"3A",X"40",X"E0",X"32",X"15",X"E5",
		X"21",X"00",X"00",X"22",X"00",X"E5",X"22",X"02",X"E5",X"C3",X"03",X"06",X"DD",X"21",X"00",X"E3",
		X"3E",X"20",X"32",X"E8",X"E0",X"DD",X"7E",X"00",X"3D",X"FA",X"00",X"02",X"21",X"0C",X"02",X"EF",
		X"11",X"10",X"00",X"DD",X"19",X"21",X"E8",X"E0",X"35",X"20",X"EA",X"C9",X"11",X"13",X"31",X"13",
		X"70",X"13",X"88",X"13",X"BC",X"13",X"C2",X"13",X"EB",X"13",X"21",X"14",X"09",X"18",X"E0",X"15",
		X"FA",X"15",X"2D",X"16",X"2D",X"16",X"49",X"16",X"5D",X"16",X"8F",X"16",X"3D",X"19",X"57",X"19",
		X"5E",X"19",X"D1",X"19",X"2F",X"1A",X"44",X"1A",X"92",X"1A",X"B9",X"1A",X"F0",X"1A",X"01",X"1B",
		X"27",X"1B",X"33",X"14",X"E0",X"18",X"AA",X"1E",X"28",X"1F",X"AC",X"20",X"C4",X"20",X"AA",X"1E",
		X"28",X"1F",X"00",X"20",X"1A",X"20",X"A4",X"1E",X"28",X"1F",X"4D",X"20",X"9C",X"20",X"23",X"1D",
		X"F3",X"1D",X"51",X"1E",X"9B",X"1E",X"9B",X"1C",X"BC",X"1C",X"14",X"1E",X"29",X"1E",X"CD",X"DC",
		X"0D",X"CD",X"0D",X"21",X"CD",X"3A",X"1B",X"CD",X"C7",X"1B",X"CD",X"A7",X"12",X"CD",X"E7",X"12",
		X"CD",X"DC",X"0D",X"3A",X"CF",X"E1",X"21",X"D0",X"E1",X"BE",X"28",X"E2",X"5F",X"16",X"E6",X"DD",
		X"21",X"00",X"00",X"DD",X"19",X"DD",X"4E",X"00",X"CB",X"21",X"20",X"11",X"21",X"CF",X"E1",X"BE",
		X"20",X"03",X"C6",X"04",X"77",X"DD",X"E5",X"C1",X"79",X"C6",X"04",X"18",X"D9",X"06",X"00",X"DD",
		X"70",X"00",X"DD",X"7E",X"01",X"21",X"A5",X"02",X"E5",X"21",X"D3",X"02",X"09",X"4E",X"23",X"66",
		X"69",X"E9",X"21",X"D0",X"E1",X"6E",X"26",X"E6",X"71",X"23",X"77",X"23",X"73",X"23",X"72",X"2C",
		X"7D",X"32",X"D0",X"E1",X"C9",X"22",X"06",X"FA",X"02",X"ED",X"02",X"22",X"03",X"2F",X"03",X"67",
		X"03",X"61",X"03",X"37",X"03",X"A6",X"0D",X"01",X"12",X"18",X"12",X"00",X"00",X"3A",X"4E",X"E0",
		X"DD",X"86",X"01",X"DD",X"77",X"01",X"DD",X"36",X"00",X"04",X"DD",X"6E",X"02",X"DD",X"66",X"03",
		X"CD",X"DB",X"03",X"7E",X"06",X"12",X"FE",X"26",X"28",X"06",X"06",X"30",X"FE",X"27",X"20",X"0D",
		X"23",X"78",X"32",X"50",X"E0",X"3A",X"50",X"E0",X"A7",X"20",X"FA",X"18",X"E6",X"CD",X"C9",X"03",
		X"18",X"E1",X"3A",X"4E",X"E0",X"DD",X"BE",X"01",X"28",X"05",X"DD",X"36",X"00",X"04",X"C9",X"DD",
		X"6E",X"02",X"DD",X"66",X"03",X"18",X"44",X"3A",X"50",X"E0",X"A7",X"20",X"0C",X"CD",X"2F",X"03",
		X"DD",X"35",X"01",X"C8",X"3E",X"04",X"32",X"50",X"E0",X"DD",X"36",X"00",X"07",X"C9",X"CD",X"DB",
		X"03",X"CD",X"C9",X"03",X"3E",X"03",X"32",X"50",X"E0",X"3A",X"50",X"E0",X"A7",X"20",X"FA",X"18",
		X"F0",X"3A",X"50",X"E0",X"A7",X"20",X"08",X"3E",X"04",X"32",X"50",X"E0",X"CD",X"FA",X"02",X"DD",
		X"36",X"00",X"08",X"C9",X"3A",X"4E",X"E0",X"CB",X"67",X"20",X"85",X"CD",X"DB",X"03",X"7E",X"23",
		X"FE",X"21",X"C8",X"FE",X"23",X"28",X"09",X"FE",X"22",X"28",X"F0",X"AF",X"12",X"13",X"18",X"EE",
		X"23",X"18",X"EB",X"7E",X"13",X"E6",X"0F",X"28",X"04",X"1B",X"CD",X"A6",X"03",X"2B",X"7E",X"1F",
		X"1F",X"1F",X"1F",X"CD",X"A7",X"03",X"7E",X"E6",X"0F",X"C6",X"30",X"12",X"13",X"C9",X"FD",X"21",
		X"00",X"04",X"FD",X"19",X"F5",X"1F",X"1F",X"1F",X"1F",X"CD",X"BD",X"03",X"F1",X"E6",X"0F",X"C6",
		X"30",X"12",X"FD",X"71",X"00",X"13",X"FD",X"23",X"C9",X"7E",X"23",X"FE",X"21",X"28",X"33",X"FE",
		X"23",X"28",X"12",X"FE",X"25",X"28",X"2D",X"FE",X"22",X"20",X"E6",X"5E",X"23",X"56",X"23",X"FD",
		X"21",X"00",X"04",X"FD",X"19",X"4E",X"23",X"3A",X"F9",X"E0",X"A7",X"C8",X"79",X"A7",X"C8",X"FE",
		X"03",X"38",X"0B",X"FE",X"06",X"28",X"03",X"FE",X"09",X"C0",X"C6",X"05",X"4F",X"C9",X"C6",X"0B",
		X"4F",X"C9",X"E1",X"C9",X"46",X"23",X"7E",X"23",X"CD",X"C1",X"03",X"10",X"FB",X"C9",X"21",X"3E",
		X"E0",X"11",X"41",X"E0",X"3A",X"00",X"D0",X"01",X"02",X"00",X"CD",X"34",X"04",X"21",X"3F",X"E0",
		X"13",X"3A",X"02",X"D0",X"1F",X"F6",X"04",X"0E",X"20",X"CD",X"34",X"04",X"3A",X"4C",X"E0",X"B0",
		X"32",X"01",X"D0",X"C9",X"1F",X"1F",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"E6",X"55",X"FE",
		X"54",X"28",X"0E",X"7E",X"E6",X"AA",X"C0",X"21",X"ED",X"E0",X"34",X"7E",X"E6",X"0F",X"C0",X"18",
		X"19",X"78",X"B1",X"47",X"3E",X"13",X"CD",X"7D",X"0D",X"1A",X"FE",X"01",X"28",X"11",X"FE",X"08",
		X"30",X"0B",X"21",X"47",X"E0",X"34",X"BE",X"C0",X"AF",X"77",X"3C",X"18",X"02",X"D6",X"08",X"21",
		X"48",X"E0",X"86",X"27",X"30",X"02",X"3E",X"99",X"77",X"C9",X"3A",X"46",X"E0",X"07",X"30",X"5B",
		X"11",X"01",X"D0",X"CB",X"67",X"28",X"07",X"3A",X"43",X"E0",X"3D",X"28",X"01",X"13",X"21",X"4A",
		X"E0",X"7E",X"23",X"77",X"2B",X"1A",X"2F",X"77",X"2B",X"E6",X"03",X"77",X"C9",X"3A",X"0B",X"E5",
		X"2A",X"F7",X"E0",X"BE",X"20",X"13",X"23",X"7E",X"54",X"5D",X"23",X"22",X"F7",X"E0",X"A7",X"28",
		X"04",X"FE",X"FF",X"20",X"D9",X"32",X"E0",X"E1",X"C9",X"21",X"4A",X"E0",X"3A",X"E0",X"E1",X"A7",
		X"28",X"13",X"3A",X"4E",X"E0",X"07",X"47",X"E6",X"01",X"3C",X"32",X"49",X"E0",X"78",X"E6",X"1E",
		X"20",X"03",X"36",X"20",X"C9",X"7E",X"36",X"FF",X"23",X"77",X"C9",X"21",X"4D",X"E0",X"3A",X"4E",
		X"E0",X"47",X"7E",X"A7",X"28",X"B7",X"FE",X"50",X"28",X"1D",X"CB",X"18",X"38",X"05",X"CB",X"18",
		X"38",X"01",X"34",X"0E",X"02",X"21",X"49",X"E0",X"FE",X"18",X"38",X"01",X"0D",X"71",X"23",X"36",
		X"00",X"FE",X"B0",X"D8",X"C3",X"7B",X"00",X"21",X"00",X"E3",X"7E",X"FE",X"04",X"20",X"0C",X"3A",
		X"09",X"E3",X"17",X"D8",X"36",X"08",X"0E",X"0A",X"C3",X"C2",X"02",X"FE",X"08",X"C8",X"21",X"4A",
		X"E0",X"36",X"20",X"23",X"36",X"00",X"C9",X"21",X"E2",X"2A",X"CD",X"00",X"03",X"3A",X"48",X"E0",
		X"C3",X"AE",X"03",X"21",X"D1",X"2A",X"CD",X"74",X"03",X"CD",X"27",X"05",X"21",X"86",X"2A",X"3A",
		X"48",X"E0",X"3D",X"28",X"03",X"21",X"97",X"2A",X"CD",X"00",X"03",X"3A",X"53",X"E0",X"E6",X"03",
		X"C8",X"1F",X"3A",X"48",X"E0",X"06",X"80",X"38",X"06",X"D6",X"01",X"27",X"C8",X"06",X"90",X"D6",
		X"01",X"27",X"F3",X"32",X"48",X"E0",X"78",X"32",X"46",X"E0",X"3C",X"FB",X"C9",X"21",X"00",X"E1",
		X"11",X"40",X"C8",X"01",X"40",X"00",X"ED",X"B0",X"1E",X"20",X"0E",X"20",X"ED",X"B0",X"1E",X"C0",
		X"0E",X"40",X"ED",X"B0",X"11",X"A0",X"C8",X"0E",X"20",X"ED",X"B0",X"0E",X"1C",X"7E",X"06",X"04",
		X"ED",X"79",X"0C",X"10",X"FB",X"23",X"3A",X"C3",X"E1",X"A7",X"28",X"2B",X"7E",X"E6",X"7F",X"01",
		X"40",X"00",X"CB",X"3F",X"30",X"01",X"04",X"20",X"F9",X"7E",X"07",X"E6",X"01",X"A8",X"5F",X"ED",
		X"A3",X"3A",X"00",X"88",X"E6",X"07",X"BB",X"C2",X"C3",X"00",X"0E",X"80",X"ED",X"A3",X"0E",X"60",
		X"ED",X"A3",X"0E",X"A0",X"ED",X"A3",X"7E",X"2F",X"D3",X"C0",X"C9",X"2A",X"DD",X"E1",X"7D",X"BC",
		X"C8",X"26",X"E0",X"7E",X"32",X"00",X"D0",X"CB",X"FF",X"32",X"00",X"D0",X"7D",X"3C",X"E6",X"07",
		X"32",X"DD",X"E1",X"C9",X"3E",X"40",X"18",X"02",X"3E",X"C0",X"32",X"50",X"E0",X"3A",X"50",X"E0",
		X"A7",X"20",X"FA",X"C9",X"21",X"00",X"E0",X"01",X"00",X"07",X"36",X"00",X"23",X"0B",X"78",X"B1",
		X"20",X"F8",X"C9",X"21",X"46",X"E0",X"7E",X"EE",X"08",X"77",X"21",X"00",X"E5",X"11",X"18",X"E5",
		X"06",X"18",X"1A",X"4F",X"7E",X"12",X"71",X"23",X"13",X"10",X"F7",X"C9",X"3A",X"46",X"E0",X"CB",
		X"5F",X"C9",X"4F",X"81",X"81",X"4F",X"06",X"00",X"21",X"0C",X"2A",X"09",X"3A",X"46",X"E0",X"A7",
		X"F0",X"11",X"00",X"E5",X"06",X"03",X"A7",X"1A",X"8E",X"27",X"12",X"13",X"23",X"10",X"F8",X"CD",
		X"AF",X"06",X"06",X"03",X"11",X"00",X"E5",X"21",X"08",X"E0",X"A7",X"1A",X"9E",X"23",X"13",X"10",
		X"FA",X"38",X"15",X"2A",X"00",X"E5",X"22",X"08",X"E0",X"3A",X"02",X"E5",X"32",X"0A",X"E0",X"3A",
		X"0E",X"E5",X"32",X"0B",X"E0",X"CD",X"85",X"06",X"11",X"84",X"80",X"CD",X"1C",X"06",X"28",X"03",
		X"11",X"A4",X"80",X"21",X"02",X"E5",X"0E",X"01",X"CD",X"E7",X"03",X"06",X"03",X"7E",X"CD",X"AE",
		X"03",X"2B",X"10",X"F9",X"C9",X"21",X"0B",X"E0",X"7E",X"0E",X"09",X"FE",X"1B",X"38",X"04",X"D6",
		X"1A",X"0E",X"06",X"C6",X"40",X"32",X"4A",X"80",X"3A",X"F9",X"E0",X"1F",X"79",X"30",X"02",X"C6",
		X"05",X"32",X"4A",X"84",X"11",X"43",X"80",X"0E",X"09",X"CD",X"E7",X"03",X"2B",X"18",X"CC",X"2A",
		X"01",X"E5",X"3A",X"45",X"E0",X"3D",X"F8",X"3D",X"28",X"01",X"24",X"CB",X"2C",X"25",X"3C",X"7C",
		X"20",X"05",X"A7",X"28",X"02",X"3E",X"FE",X"21",X"03",X"E5",X"BE",X"C0",X"7E",X"FE",X"03",X"C8",
		X"34",X"21",X"15",X"E5",X"34",X"3A",X"15",X"E5",X"3D",X"28",X"03",X"4F",X"3E",X"01",X"21",X"7C",
		X"80",X"CD",X"EC",X"06",X"CD",X"EC",X"06",X"28",X"03",X"79",X"C6",X"30",X"77",X"23",X"A7",X"C8",
		X"3C",X"C9",X"21",X"40",X"E0",X"3A",X"03",X"D0",X"47",X"3C",X"E6",X"03",X"20",X"02",X"3E",X"05",
		X"77",X"23",X"78",X"0F",X"0F",X"47",X"E6",X"03",X"32",X"45",X"E0",X"3A",X"04",X"D0",X"CB",X"57",
		X"78",X"28",X"1F",X"1F",X"1F",X"ED",X"44",X"E6",X"0F",X"CB",X"5F",X"28",X"01",X"3C",X"77",X"23",
		X"77",X"3A",X"04",X"D0",X"2F",X"1F",X"47",X"E6",X"01",X"23",X"77",X"78",X"1F",X"E6",X"01",X"23",
		X"77",X"C9",X"1F",X"1F",X"2F",X"47",X"3C",X"E6",X"03",X"77",X"78",X"1F",X"1F",X"E6",X"03",X"FE",
		X"02",X"DE",X"F5",X"18",X"DA",X"CD",X"29",X"0D",X"21",X"97",X"2C",X"CD",X"00",X"03",X"CD",X"27",
		X"05",X"21",X"57",X"2C",X"CD",X"4E",X"03",X"11",X"54",X"E0",X"01",X"20",X"00",X"3A",X"44",X"E0",
		X"A7",X"20",X"34",X"CD",X"9F",X"07",X"CD",X"E8",X"07",X"7E",X"FE",X"32",X"20",X"20",X"3E",X"53",
		X"32",X"5F",X"E0",X"32",X"68",X"E0",X"21",X"62",X"E0",X"7E",X"87",X"D6",X"30",X"FE",X"3A",X"38",
		X"06",X"D6",X"0A",X"77",X"2B",X"3E",X"31",X"77",X"21",X"54",X"E0",X"CD",X"4E",X"03",X"3A",X"47",
		X"E0",X"A7",X"20",X"FA",X"C3",X"E8",X"05",X"CD",X"D3",X"07",X"CD",X"DD",X"07",X"18",X"E9",X"21",
		X"67",X"2C",X"ED",X"B0",X"21",X"57",X"E0",X"3A",X"41",X"E0",X"11",X"08",X"00",X"FE",X"08",X"38",
		X"12",X"C6",X"28",X"77",X"19",X"36",X"53",X"23",X"23",X"23",X"36",X"31",X"11",X"06",X"00",X"19",
		X"36",X"00",X"C9",X"3D",X"C8",X"11",X"0B",X"00",X"19",X"C6",X"31",X"77",X"11",X"06",X"00",X"19",
		X"36",X"53",X"C9",X"21",X"7D",X"2C",X"ED",X"B0",X"21",X"5B",X"E0",X"18",X"CA",X"CD",X"E8",X"07",
		X"21",X"5B",X"E0",X"3A",X"42",X"E0",X"18",X"C2",X"21",X"54",X"E0",X"CD",X"4E",X"03",X"2A",X"54",
		X"E0",X"11",X"40",X"00",X"19",X"22",X"54",X"E0",X"21",X"57",X"E0",X"34",X"C9",X"21",X"77",X"E2",
		X"06",X"07",X"7E",X"A7",X"28",X"0B",X"2B",X"10",X"F9",X"C9",X"21",X"61",X"E2",X"06",X"12",X"18",
		X"F1",X"34",X"7D",X"D6",X"50",X"87",X"87",X"DD",X"77",X"01",X"C9",X"DD",X"7E",X"07",X"E6",X"F8",
		X"6F",X"26",X"20",X"29",X"29",X"DD",X"7E",X"03",X"1F",X"57",X"1F",X"1F",X"E6",X"1F",X"85",X"6F",
		X"C9",X"3A",X"00",X"E3",X"FE",X"06",X"30",X"7A",X"3A",X"E2",X"E1",X"DD",X"96",X"0F",X"ED",X"44",
		X"DD",X"77",X"03",X"FE",X"E0",X"38",X"6D",X"DD",X"4E",X"0B",X"0D",X"20",X"6B",X"FE",X"E8",X"30",
		X"67",X"E1",X"DD",X"36",X"00",X"00",X"DD",X"7E",X"0D",X"37",X"17",X"D8",X"37",X"17",X"21",X"18",
		X"2E",X"30",X"01",X"24",X"5F",X"16",X"00",X"19",X"46",X"DD",X"5E",X"01",X"16",X"E1",X"78",X"17",
		X"30",X"10",X"06",X"01",X"17",X"38",X"27",X"7B",X"FE",X"60",X"38",X"06",X"62",X"D6",X"5E",X"6F",
		X"36",X"00",X"FD",X"21",X"00",X"00",X"FD",X"19",X"7B",X"1F",X"1F",X"E6",X"3F",X"C6",X"50",X"6F",
		X"26",X"E2",X"11",X"04",X"00",X"FD",X"72",X"02",X"FD",X"19",X"10",X"F9",X"72",X"C9",X"CD",X"82",
		X"08",X"21",X"74",X"E1",X"01",X"00",X"18",X"71",X"23",X"10",X"FC",X"21",X"D1",X"E1",X"70",X"23",
		X"70",X"C9",X"E1",X"C9",X"DD",X"36",X"0B",X"01",X"DD",X"7E",X"0D",X"07",X"D8",X"17",X"21",X"18",
		X"2E",X"30",X"01",X"24",X"5F",X"16",X"00",X"19",X"DD",X"5E",X"01",X"16",X"E1",X"FD",X"21",X"00",
		X"00",X"FD",X"19",X"56",X"23",X"5E",X"23",X"4E",X"06",X"00",X"21",X"F5",X"08",X"09",X"4E",X"23",
		X"66",X"69",X"DD",X"4E",X"03",X"DD",X"7E",X"07",X"CD",X"ED",X"08",X"AF",X"E9",X"2F",X"47",X"3A",
		X"3C",X"E0",X"80",X"47",X"C9",X"69",X"09",X"5A",X"09",X"CF",X"09",X"CD",X"09",X"F5",X"0A",X"43",
		X"09",X"E2",X"0A",X"90",X"0A",X"56",X"0A",X"B7",X"0A",X"52",X"0A",X"9F",X"0A",X"C9",X"09",X"25",
		X"0B",X"76",X"09",X"97",X"09",X"BA",X"09",X"1E",X"0A",X"44",X"0A",X"34",X"09",X"25",X"09",X"1D",
		X"0B",X"B0",X"09",X"83",X"09",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"E6",X"1F",X"FE",X"0B",X"38",
		X"38",X"1C",X"18",X"35",X"3A",X"4E",X"E0",X"E6",X"03",X"28",X"01",X"14",X"CD",X"69",X"09",X"16",
		X"3B",X"18",X"1B",X"FD",X"21",X"A4",X"E1",X"FD",X"77",X"0A",X"FD",X"77",X"0E",X"FD",X"77",X"12",
		X"FD",X"77",X"16",X"CD",X"95",X"0A",X"3E",X"F8",X"80",X"47",X"CD",X"69",X"09",X"14",X"3E",X"10",
		X"81",X"4F",X"21",X"04",X"00",X"EB",X"FD",X"19",X"EB",X"DD",X"7E",X"0B",X"A7",X"79",X"20",X"35",
		X"C6",X"08",X"FE",X"20",X"38",X"35",X"FD",X"70",X"00",X"FD",X"73",X"01",X"FD",X"72",X"02",X"FD",
		X"71",X"03",X"C9",X"DD",X"7E",X"08",X"1E",X"07",X"CB",X"3F",X"CB",X"13",X"C6",X"7A",X"57",X"78",
		X"FE",X"80",X"D2",X"25",X"0B",X"18",X"DF",X"3E",X"08",X"80",X"47",X"FD",X"21",X"74",X"E1",X"79",
		X"FE",X"F8",X"D0",X"18",X"D1",X"C6",X"08",X"FE",X"F0",X"38",X"CB",X"FD",X"36",X"02",X"00",X"C9",
		X"3A",X"4E",X"E0",X"CB",X"57",X"28",X"BF",X"14",X"18",X"BC",X"3E",X"0E",X"80",X"60",X"47",X"2E",
		X"01",X"CD",X"E4",X"09",X"11",X"08",X"76",X"18",X"11",X"3E",X"0A",X"18",X"02",X"3E",X"05",X"80",
		X"60",X"47",X"2E",X"01",X"CD",X"E4",X"09",X"11",X"08",X"71",X"44",X"21",X"08",X"00",X"EB",X"FD",
		X"19",X"EB",X"2E",X"00",X"CD",X"69",X"09",X"FD",X"70",X"04",X"2D",X"20",X"29",X"3E",X"40",X"AB",
		X"FD",X"77",X"05",X"3E",X"08",X"FD",X"72",X"06",X"81",X"FD",X"77",X"07",X"C6",X"08",X"FE",X"F8",
		X"30",X"0A",X"FE",X"20",X"D0",X"DD",X"7E",X"0B",X"A7",X"28",X"06",X"C9",X"DD",X"7E",X"0B",X"A7",
		X"C8",X"FD",X"36",X"06",X"00",X"C9",X"14",X"FD",X"73",X"05",X"3E",X"10",X"18",X"D7",X"C5",X"D5",
		X"21",X"02",X"08",X"09",X"44",X"4D",X"79",X"C6",X"08",X"FE",X"D0",X"30",X"11",X"CD",X"83",X"09",
		X"11",X"04",X"00",X"FD",X"19",X"D1",X"C1",X"2E",X"00",X"FD",X"75",X"0A",X"18",X"A6",X"FD",X"36",
		X"02",X"00",X"18",X"EC",X"32",X"A6",X"E1",X"32",X"AA",X"E1",X"32",X"AE",X"E1",X"CD",X"95",X"0A",
		X"18",X"10",X"3E",X"18",X"18",X"02",X"3E",X"0D",X"FD",X"21",X"74",X"E1",X"80",X"47",X"3E",X"F8",
		X"81",X"4F",X"AF",X"CD",X"6F",X"0A",X"EB",X"11",X"08",X"00",X"FD",X"19",X"EB",X"3E",X"10",X"81",
		X"6F",X"FD",X"77",X"03",X"FD",X"77",X"07",X"FD",X"70",X"00",X"3E",X"F0",X"80",X"FD",X"77",X"04",
		X"FD",X"73",X"01",X"FD",X"73",X"05",X"FD",X"72",X"02",X"14",X"14",X"FD",X"72",X"06",X"15",X"C9",
		X"CD",X"95",X"0A",X"18",X"CD",X"3A",X"F9",X"E0",X"1F",X"D0",X"7B",X"F6",X"0C",X"5F",X"C9",X"FD",
		X"21",X"74",X"E1",X"FD",X"36",X"0A",X"00",X"FD",X"36",X"0E",X"00",X"3E",X"18",X"80",X"47",X"AF",
		X"CD",X"6F",X"0A",X"FD",X"72",X"06",X"C9",X"3E",X"18",X"80",X"47",X"FD",X"21",X"74",X"E1",X"3E",
		X"F8",X"CD",X"CD",X"0A",X"21",X"0C",X"00",X"EB",X"FD",X"19",X"EB",X"3E",X"08",X"CD",X"6F",X"0A",
		X"FD",X"75",X"0B",X"D6",X"10",X"FD",X"77",X"08",X"FD",X"77",X"09",X"7A",X"C6",X"03",X"FD",X"77",
		X"0A",X"C9",X"FD",X"21",X"A4",X"E1",X"FD",X"77",X"06",X"CD",X"95",X"0A",X"21",X"08",X"F8",X"09",
		X"44",X"4D",X"C3",X"76",X"09",X"FD",X"21",X"A4",X"E1",X"FD",X"36",X"1A",X"00",X"CD",X"95",X"0A",
		X"3E",X"F8",X"CD",X"13",X"0B",X"3E",X"08",X"CD",X"0C",X"0B",X"3E",X"18",X"EB",X"11",X"08",X"00",
		X"FD",X"19",X"EB",X"CD",X"6F",X"0A",X"7A",X"C6",X"02",X"FD",X"77",X"06",X"C9",X"3A",X"4E",X"E0",
		X"CB",X"4F",X"28",X"01",X"1C",X"CD",X"76",X"09",X"DD",X"7E",X"01",X"FE",X"60",X"D8",X"EB",X"11",
		X"A0",X"FF",X"FD",X"19",X"EB",X"C3",X"76",X"09",X"CD",X"8E",X"0C",X"CD",X"BF",X"0C",X"3A",X"04",
		X"D0",X"CB",X"6F",X"C0",X"21",X"A9",X"2A",X"CD",X"00",X"03",X"3E",X"FF",X"32",X"51",X"E0",X"21",
		X"53",X"E0",X"7E",X"4E",X"A9",X"A1",X"1F",X"38",X"08",X"3A",X"51",X"E0",X"47",X"79",X"10",X"F3",
		X"C9",X"21",X"0E",X"E5",X"7E",X"3C",X"FE",X"34",X"30",X"E0",X"77",X"2A",X"16",X"E5",X"46",X"23",
		X"7E",X"E6",X"7F",X"23",X"FE",X"06",X"20",X"F6",X"78",X"32",X"0B",X"E5",X"22",X"16",X"E5",X"32",
		X"23",X"E5",X"22",X"2E",X"E5",X"CD",X"12",X"0D",X"18",X"C0",X"CD",X"B1",X"0C",X"21",X"94",X"26",
		X"22",X"16",X"E5",X"C3",X"BF",X"0C",X"2A",X"16",X"E5",X"2B",X"7E",X"2B",X"E6",X"7F",X"FE",X"06",
		X"20",X"F7",X"11",X"DC",X"E1",X"EB",X"7E",X"36",X"00",X"EB",X"A7",X"20",X"EC",X"7E",X"32",X"0B",
		X"E5",X"23",X"23",X"22",X"16",X"E5",X"C9",X"21",X"00",X"E1",X"01",X"00",X"04",X"CD",X"FA",X"05",
		X"DD",X"21",X"00",X"E3",X"DD",X"36",X"00",X"01",X"DD",X"36",X"10",X"09",X"DD",X"36",X"01",X"B0",
		X"DD",X"36",X"21",X"A0",X"DD",X"21",X"70",X"E3",X"3E",X"60",X"06",X"09",X"11",X"10",X"00",X"DD",
		X"77",X"01",X"DD",X"19",X"C6",X"04",X"10",X"F7",X"CD",X"96",X"0B",X"2B",X"46",X"3E",X"04",X"21",
		X"00",X"C0",X"05",X"F2",X"FA",X"0B",X"3E",X"07",X"26",X"A8",X"32",X"14",X"E5",X"22",X"06",X"E3",
		X"3E",X"02",X"32",X"08",X"E5",X"CD",X"8D",X"0D",X"3A",X"13",X"E5",X"3D",X"FE",X"05",X"CE",X"00",
		X"06",X"FB",X"1F",X"38",X"01",X"04",X"78",X"32",X"C5",X"E1",X"CD",X"81",X"29",X"A7",X"20",X"5F",
		X"21",X"0F",X"E5",X"CB",X"46",X"20",X"58",X"34",X"3A",X"10",X"E5",X"A7",X"28",X"58",X"21",X"5F",
		X"2A",X"CD",X"00",X"03",X"3A",X"10",X"E5",X"FE",X"04",X"38",X"02",X"3E",X"03",X"C6",X"30",X"32",
		X"56",X"81",X"3E",X"1C",X"CD",X"6F",X"0D",X"3E",X"40",X"32",X"0A",X"E3",X"0E",X"68",X"21",X"B6",
		X"30",X"46",X"CB",X"78",X"20",X"14",X"23",X"5E",X"23",X"7E",X"23",X"EB",X"26",X"83",X"71",X"26",
		X"87",X"70",X"0C",X"2C",X"BD",X"20",X"F5",X"EB",X"18",X"E7",X"3E",X"D3",X"21",X"D8",X"30",X"11",
		X"10",X"E2",X"46",X"CB",X"78",X"20",X"08",X"12",X"13",X"10",X"FC",X"3C",X"23",X"18",X"F3",X"21",
		X"46",X"E0",X"34",X"C3",X"6E",X"02",X"21",X"47",X"2A",X"CD",X"00",X"03",X"18",X"B4",X"AF",X"32",
		X"4D",X"E0",X"CD",X"95",X"0C",X"CD",X"03",X"06",X"21",X"00",X"E5",X"01",X"16",X"00",X"CD",X"FA",
		X"05",X"32",X"0F",X"E5",X"3A",X"40",X"E0",X"32",X"15",X"E5",X"21",X"62",X"21",X"22",X"16",X"E5",
		X"C9",X"21",X"DE",X"26",X"22",X"F7",X"E0",X"21",X"03",X"E5",X"01",X"11",X"00",X"18",X"DF",X"CD",
		X"29",X"0D",X"21",X"21",X"84",X"0E",X"06",X"3A",X"0E",X"E5",X"FE",X"1A",X"3E",X"00",X"38",X"01",
		X"3C",X"32",X"F9",X"E0",X"C5",X"0E",X"01",X"CD",X"E7",X"03",X"79",X"C1",X"06",X"1E",X"77",X"23",
		X"10",X"FC",X"23",X"23",X"0D",X"20",X"F5",X"21",X"0F",X"2B",X"CD",X"00",X"03",X"CD",X"68",X"06",
		X"CD",X"85",X"06",X"3A",X"46",X"E0",X"CB",X"67",X"28",X"0F",X"CD",X"03",X"06",X"CD",X"68",X"06",
		X"CD",X"03",X"06",X"21",X"72",X"2B",X"CD",X"00",X"03",X"CD",X"D5",X"06",X"CD",X"2C",X"21",X"CD",
		X"8A",X"29",X"3A",X"0E",X"E5",X"0E",X"02",X"FE",X"1A",X"38",X"04",X"D6",X"1A",X"0E",X"07",X"C6",
		X"40",X"32",X"52",X"80",X"79",X"32",X"52",X"84",X"C9",X"21",X"00",X"80",X"01",X"00",X"08",X"CD",
		X"FA",X"05",X"21",X"00",X"E1",X"01",X"C6",X"00",X"CD",X"FA",X"05",X"3A",X"43",X"E0",X"3D",X"28",
		X"09",X"21",X"46",X"E0",X"AF",X"CB",X"5E",X"28",X"01",X"3C",X"32",X"4C",X"E0",X"21",X"04",X"D0",
		X"AE",X"21",X"3C",X"E0",X"36",X"EF",X"16",X"FF",X"1F",X"30",X"03",X"14",X"36",X"F1",X"23",X"72",
		X"01",X"00",X"40",X"AF",X"ED",X"79",X"0C",X"10",X"FB",X"F3",X"CD",X"7D",X"0D",X"FB",X"C9",X"F3",
		X"CD",X"75",X"0D",X"FB",X"C9",X"E5",X"21",X"46",X"E0",X"CB",X"7E",X"E1",X"F0",X"E5",X"2A",X"DE",
		X"E1",X"26",X"E0",X"77",X"7D",X"3C",X"E6",X"07",X"32",X"DE",X"E1",X"E1",X"C9",X"CD",X"48",X"29",
		X"CD",X"C2",X"0C",X"06",X"20",X"C5",X"CD",X"06",X"11",X"21",X"E2",X"E1",X"7E",X"C6",X"08",X"77",
		X"C1",X"10",X"F2",X"C3",X"3B",X"0D",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"01",X"4A",X"30",X"81",
		X"4F",X"0A",X"4F",X"EB",X"11",X"20",X"00",X"7E",X"A7",X"20",X"03",X"19",X"18",X"F9",X"22",X"54",
		X"E0",X"0A",X"03",X"3D",X"C8",X"F2",X"CD",X"0D",X"3C",X"77",X"19",X"18",X"F4",X"3A",X"54",X"E0",
		X"3C",X"6F",X"E6",X"1F",X"20",X"E8",X"7D",X"D6",X"20",X"6F",X"18",X"E2",X"CD",X"5B",X"12",X"3A",
		X"E2",X"E1",X"21",X"09",X"E5",X"47",X"AE",X"E6",X"F8",X"C8",X"78",X"E6",X"F8",X"77",X"CD",X"06",
		X"11",X"3A",X"4D",X"E0",X"A7",X"C0",X"21",X"0B",X"E5",X"34",X"7E",X"5F",X"A7",X"28",X"07",X"E6",
		X"1F",X"20",X"03",X"CD",X"D6",X"29",X"7B",X"2A",X"16",X"E5",X"BE",X"20",X"0B",X"23",X"7E",X"E6",
		X"7F",X"32",X"D7",X"E1",X"23",X"22",X"16",X"E5",X"21",X"D7",X"E1",X"7E",X"3D",X"F8",X"36",X"00",
		X"FE",X"18",X"D2",X"45",X"0F",X"FE",X"17",X"28",X"26",X"D6",X"06",X"FA",X"8A",X"0E",X"D6",X"07",
		X"FA",X"F0",X"0E",X"87",X"87",X"87",X"5F",X"16",X"00",X"FD",X"21",X"00",X"10",X"FD",X"19",X"CD",
		X"93",X"0E",X"FD",X"7E",X"06",X"A7",X"28",X"03",X"CD",X"FD",X"07",X"DD",X"71",X"00",X"C9",X"3E",
		X"19",X"32",X"70",X"E3",X"C9",X"3E",X"01",X"32",X"DC",X"E1",X"2A",X"E4",X"E0",X"7D",X"E6",X"1F",
		X"F6",X"C0",X"6F",X"36",X"0A",X"01",X"20",X"00",X"5D",X"09",X"36",X"0B",X"7B",X"3D",X"E6",X"1F",
		X"F6",X"C0",X"6F",X"CD",X"81",X"29",X"C6",X"41",X"77",X"22",X"DA",X"E1",X"09",X"36",X"F2",X"01",
		X"E0",X"03",X"09",X"3A",X"F9",X"E0",X"C6",X"05",X"77",X"C9",X"3C",X"28",X"C8",X"C6",X"05",X"32",
		X"08",X"E5",X"C9",X"FD",X"7E",X"00",X"FE",X"02",X"28",X"1B",X"FE",X"07",X"38",X"1C",X"16",X"00",
		X"FD",X"5E",X"05",X"DD",X"21",X"70",X"E3",X"FD",X"46",X"04",X"DD",X"7E",X"00",X"A7",X"28",X"13",
		X"DD",X"19",X"10",X"F6",X"C9",X"21",X"D7",X"E1",X"36",X"11",X"11",X"F0",X"FF",X"DD",X"21",X"F0",
		X"E4",X"18",X"E4",X"FD",X"7E",X"00",X"DD",X"77",X"0C",X"FD",X"7E",X"01",X"DD",X"77",X"0D",X"3A",
		X"09",X"E5",X"D6",X"02",X"DD",X"77",X"0F",X"CD",X"3D",X"15",X"FD",X"86",X"03",X"DD",X"77",X"07",
		X"DD",X"36",X"0B",X"00",X"DD",X"36",X"03",X"00",X"DD",X"36",X"0E",X"00",X"FD",X"4E",X"02",X"C9",
		X"3C",X"CA",X"40",X"0F",X"F5",X"FD",X"21",X"4E",X"10",X"CD",X"BA",X"0E",X"F1",X"C6",X"86",X"DD",
		X"77",X"0D",X"DD",X"71",X"00",X"21",X"4A",X"30",X"85",X"C6",X"80",X"6F",X"6E",X"FD",X"2A",X"E4",
		X"E0",X"11",X"20",X"00",X"7E",X"23",X"3D",X"F2",X"22",X"0F",X"3C",X"FD",X"77",X"00",X"FD",X"19",
		X"18",X"F2",X"C8",X"22",X"E6",X"E0",X"3D",X"28",X"11",X"FD",X"21",X"55",X"10",X"CD",X"9E",X"0E",
		X"DD",X"36",X"0A",X"00",X"DD",X"34",X"0E",X"DD",X"71",X"00",X"3E",X"0D",X"32",X"D7",X"E1",X"C9",
		X"2A",X"E6",X"E0",X"18",X"C8",X"D6",X"1F",X"FA",X"B7",X"0F",X"21",X"C5",X"E1",X"0E",X"FF",X"23",
		X"0C",X"D6",X"08",X"F2",X"4F",X"0F",X"C6",X"08",X"28",X"10",X"77",X"23",X"23",X"23",X"77",X"23",
		X"23",X"23",X"77",X"0D",X"F8",X"21",X"D6",X"E1",X"34",X"C9",X"77",X"FD",X"21",X"70",X"E3",X"11",
		X"10",X"00",X"06",X"19",X"0D",X"FA",X"A5",X"0F",X"FD",X"7E",X"00",X"D6",X"22",X"FE",X"06",X"30",
		X"19",X"6F",X"CB",X"4D",X"20",X"14",X"61",X"FD",X"7E",X"0D",X"FE",X"2A",X"20",X"01",X"24",X"25",
		X"20",X"08",X"CB",X"55",X"20",X"09",X"FD",X"36",X"00",X"24",X"FD",X"19",X"10",X"DA",X"C9",X"FD",
		X"36",X"0F",X"01",X"18",X"F5",X"FD",X"7E",X"00",X"D6",X"1E",X"FE",X"02",X"30",X"04",X"FD",X"36",
		X"00",X"24",X"FD",X"19",X"10",X"EF",X"C9",X"C6",X"08",X"FE",X"04",X"30",X"08",X"21",X"0B",X"E5",
		X"46",X"23",X"70",X"23",X"77",X"3A",X"D5",X"E1",X"A7",X"C8",X"5F",X"16",X"00",X"FD",X"21",X"FF",
		X"E3",X"FD",X"19",X"21",X"70",X"E3",X"1E",X"10",X"01",X"3A",X"05",X"7E",X"A7",X"CA",X"5D",X"10",
		X"19",X"10",X"F8",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A5",
		X"00",X"0E",X"12",X"F0",X"10",X"00",X"01",X"00",X"01",X"0F",X"12",X"F0",X"10",X"00",X"01",X"00",
		X"02",X"10",X"12",X"F0",X"10",X"00",X"01",X"00",X"03",X"11",X"12",X"F0",X"10",X"00",X"01",X"00",
		X"0D",X"25",X"12",X"FD",X"06",X"10",X"00",X"00",X"0A",X"21",X"1D",X"F0",X"05",X"10",X"00",X"00",
		X"04",X"12",X"16",X"F4",X"18",X"10",X"01",X"00",X"05",X"16",X"16",X"F2",X"18",X"10",X"01",X"00",
		X"06",X"1B",X"16",X"F0",X"18",X"10",X"01",X"00",X"0B",X"23",X"17",X"F0",X"01",X"20",X"00",X"00",
		X"13",X"00",X"10",X"00",X"00",X"00",X"4A",X"14",X"00",X"03",X"40",X"00",X"00",X"EB",X"DD",X"21",
		X"00",X"00",X"DD",X"19",X"DD",X"71",X"0D",X"DD",X"36",X"09",X"00",X"DD",X"36",X"08",X"00",X"FD",
		X"56",X"07",X"DD",X"72",X"07",X"FD",X"7E",X"00",X"D6",X"1E",X"FE",X"0A",X"D0",X"CB",X"4F",X"C0",
		X"FD",X"7E",X"03",X"D6",X"10",X"FE",X"E0",X"D0",X"79",X"FE",X"3A",X"28",X"36",X"CD",X"92",X"20",
		X"ED",X"5F",X"E6",X"7F",X"47",X"3A",X"03",X"E3",X"80",X"D6",X"2F",X"4F",X"DD",X"96",X"03",X"C6",
		X"08",X"FE",X"11",X"79",X"30",X"03",X"EE",X"10",X"4F",X"FD",X"BE",X"03",X"17",X"DD",X"77",X"0C",
		X"79",X"CD",X"38",X"15",X"92",X"1F",X"1F",X"1F",X"E6",X"1F",X"C6",X"02",X"41",X"CB",X"38",X"0E",
		X"2E",X"18",X"0F",X"01",X"2A",X"8F",X"CB",X"3A",X"CB",X"3A",X"CB",X"3A",X"3A",X"14",X"E5",X"EE",
		X"1F",X"92",X"21",X"00",X"31",X"85",X"6F",X"56",X"FD",X"7E",X"03",X"DD",X"77",X"03",X"CB",X"3F",
		X"90",X"30",X"02",X"ED",X"44",X"1E",X"FF",X"1C",X"92",X"30",X"FC",X"82",X"DD",X"73",X"05",X"06",
		X"08",X"CB",X"27",X"BA",X"CB",X"13",X"CB",X"43",X"20",X"01",X"92",X"10",X"F4",X"7B",X"2F",X"DD",
		X"77",X"04",X"DD",X"71",X"00",X"C9",X"21",X"D9",X"E1",X"7E",X"A7",X"C2",X"9A",X"11",X"3A",X"08",
		X"E5",X"FE",X"03",X"30",X"79",X"47",X"05",X"21",X"B4",X"2C",X"3A",X"E2",X"E1",X"1F",X"1F",X"1F",
		X"E6",X"1F",X"85",X"10",X"02",X"C6",X"20",X"6F",X"4E",X"3A",X"E2",X"E1",X"1F",X"1F",X"1F",X"E6",
		X"1F",X"5F",X"16",X"83",X"FD",X"21",X"00",X"04",X"FD",X"19",X"EB",X"11",X"20",X"00",X"06",X"07",
		X"3A",X"14",X"E5",X"B8",X"28",X"07",X"36",X"00",X"19",X"FD",X"19",X"10",X"F6",X"22",X"E4",X"E0",
		X"71",X"FD",X"36",X"00",X"04",X"19",X"FD",X"19",X"36",X"F3",X"FD",X"36",X"00",X"04",X"10",X"F5",
		X"3A",X"E2",X"E1",X"1F",X"1F",X"E6",X"3E",X"C6",X"00",X"6F",X"26",X"E2",X"3A",X"14",X"E5",X"EE",
		X"1F",X"57",X"FD",X"21",X"24",X"2C",X"FD",X"09",X"FD",X"7E",X"00",X"5F",X"E6",X"70",X"07",X"B2",
		X"07",X"07",X"07",X"77",X"E6",X"F8",X"57",X"7B",X"E6",X"07",X"B2",X"23",X"77",X"C9",X"87",X"C6",
		X"7A",X"77",X"87",X"28",X"02",X"3E",X"0A",X"32",X"D8",X"E1",X"4E",X"CB",X"19",X"D8",X"CB",X"19",
		X"21",X"D8",X"E1",X"35",X"F2",X"B6",X"11",X"36",X"0B",X"3A",X"14",X"E5",X"38",X"3C",X"FE",X"07",
		X"28",X"3E",X"3E",X"0B",X"18",X"27",X"7E",X"21",X"14",X"E5",X"30",X"1C",X"A7",X"20",X"01",X"35",
		X"C6",X"F3",X"FE",X"FC",X"38",X"02",X"D6",X"0C",X"4F",X"C6",X"03",X"FA",X"C9",X"11",X"C2",X"29",
		X"11",X"79",X"D6",X"10",X"4F",X"C3",X"29",X"11",X"FE",X"09",X"20",X"01",X"34",X"2F",X"C6",X"F2",
		X"FE",X"F0",X"30",X"02",X"C6",X"0C",X"4F",X"C3",X"29",X"11",X"FE",X"04",X"3E",X"0B",X"20",X"D0",
		X"21",X"D9",X"E1",X"34",X"2A",X"E1",X"E1",X"22",X"F1",X"E0",X"21",X"00",X"00",X"22",X"EF",X"E0",
		X"C9",X"21",X"44",X"2D",X"ED",X"53",X"EB",X"E0",X"22",X"E9",X"E0",X"3A",X"4E",X"E0",X"C6",X"03",
		X"DD",X"77",X"01",X"DD",X"36",X"00",X"0B",X"C9",X"3A",X"4E",X"E0",X"DD",X"BE",X"01",X"20",X"F3",
		X"2A",X"EB",X"E0",X"23",X"22",X"EB",X"E0",X"2B",X"EB",X"FD",X"21",X"00",X"04",X"FD",X"19",X"2A",
		X"E9",X"E0",X"01",X"20",X"00",X"7E",X"23",X"3D",X"FE",X"03",X"38",X"0D",X"3C",X"12",X"FD",X"36",
		X"00",X"80",X"EB",X"09",X"EB",X"FD",X"09",X"18",X"EC",X"3D",X"FA",X"55",X"12",X"28",X"B9",X"5E",
		X"23",X"56",X"23",X"18",X"AF",X"21",X"97",X"2C",X"C3",X"00",X"03",X"3A",X"0D",X"E5",X"3D",X"F8",
		X"21",X"AB",X"2C",X"3A",X"4E",X"E0",X"E6",X"3F",X"28",X"1B",X"E6",X"1F",X"C0",X"CD",X"7B",X"03",
		X"CD",X"88",X"12",X"36",X"02",X"EB",X"36",X"12",X"21",X"0B",X"E5",X"7E",X"23",X"96",X"FE",X"40",
		X"D8",X"23",X"36",X"00",X"C9",X"CD",X"00",X"03",X"3A",X"0D",X"E5",X"21",X"55",X"80",X"01",X"02",
		X"13",X"11",X"20",X"00",X"3D",X"28",X"08",X"19",X"0C",X"05",X"3D",X"28",X"02",X"04",X"19",X"70",
		X"11",X"00",X"04",X"EB",X"19",X"71",X"C9",X"21",X"70",X"E3",X"11",X"10",X"00",X"01",X"02",X"19",
		X"7E",X"FE",X"14",X"28",X"2A",X"FE",X"1E",X"38",X"1B",X"FE",X"20",X"38",X"08",X"FE",X"22",X"38",
		X"13",X"FE",X"2A",X"30",X"0F",X"3A",X"DF",X"E1",X"1F",X"1F",X"D8",X"79",X"32",X"DF",X"E1",X"C6",
		X"15",X"C3",X"6F",X"0D",X"19",X"10",X"D9",X"3A",X"DF",X"E1",X"A7",X"C8",X"AF",X"18",X"ED",X"3A",
		X"DF",X"E1",X"1F",X"0D",X"30",X"E5",X"C9",X"3A",X"DC",X"E1",X"A7",X"C8",X"3A",X"4E",X"E0",X"E6",
		X"0F",X"28",X"04",X"E6",X"07",X"C0",X"3C",X"3C",X"4F",X"2A",X"DA",X"E1",X"7E",X"D6",X"5A",X"28",
		X"0A",X"3C",X"06",X"04",X"C6",X"05",X"28",X"03",X"10",X"FA",X"C9",X"11",X"00",X"04",X"19",X"71",
		X"C9",X"21",X"00",X"40",X"22",X"02",X"E3",X"3A",X"4E",X"E0",X"E6",X"03",X"20",X"48",X"DD",X"35",
		X"0A",X"F2",X"66",X"13",X"21",X"5F",X"2A",X"CD",X"7B",X"03",X"3E",X"18",X"CD",X"75",X"0D",X"18",
		X"29",X"CD",X"48",X"15",X"07",X"07",X"30",X"2B",X"2A",X"1A",X"E3",X"11",X"79",X"FF",X"19",X"7C",
		X"A7",X"20",X"05",X"7D",X"FE",X"D1",X"38",X"02",X"3E",X"D1",X"5F",X"CB",X"3B",X"83",X"2F",X"6F",
		X"3E",X"FF",X"DE",X"00",X"67",X"2B",X"67",X"22",X"08",X"E3",X"DD",X"34",X"00",X"CD",X"76",X"15",
		X"C3",X"B8",X"08",X"CD",X"8A",X"14",X"CD",X"33",X"15",X"D6",X"1C",X"32",X"07",X"E3",X"18",X"ED",
		X"DD",X"34",X"00",X"3E",X"14",X"CD",X"75",X"0D",X"CD",X"48",X"15",X"2A",X"0E",X"E3",X"CD",X"A4",
		X"14",X"CD",X"33",X"15",X"D6",X"1E",X"18",X"E3",X"CD",X"48",X"15",X"2A",X"0E",X"E3",X"CD",X"A4",
		X"14",X"2A",X"06",X"E3",X"ED",X"5B",X"08",X"E3",X"19",X"22",X"06",X"E3",X"21",X"0C",X"00",X"19",
		X"22",X"08",X"E3",X"CB",X"14",X"38",X"0F",X"CD",X"33",X"15",X"D6",X"1D",X"47",X"3A",X"07",X"E3",
		X"B8",X"38",X"03",X"DD",X"34",X"00",X"CD",X"AC",X"15",X"C3",X"B8",X"08",X"DD",X"36",X"00",X"02",
		X"18",X"B6",X"2A",X"02",X"E3",X"ED",X"5B",X"04",X"E3",X"19",X"22",X"02",X"E3",X"2A",X"06",X"E3",
		X"ED",X"5B",X"08",X"E3",X"19",X"22",X"06",X"E3",X"CD",X"B8",X"08",X"DD",X"35",X"0A",X"C0",X"DD",
		X"34",X"00",X"DD",X"36",X"0D",X"03",X"3E",X"1F",X"C3",X"75",X"0D",X"AF",X"32",X"A2",X"E1",X"DD",
		X"35",X"0A",X"F0",X"DD",X"7E",X"0D",X"FE",X"09",X"D2",X"18",X"01",X"FE",X"05",X"38",X"0B",X"CD",
		X"B8",X"08",X"DD",X"34",X"0D",X"DD",X"36",X"0A",X"0E",X"C9",X"DD",X"CB",X"0A",X"4E",X"C0",X"EE",
		X"07",X"DD",X"77",X"0D",X"DD",X"7E",X"0A",X"FE",X"C0",X"D2",X"B8",X"08",X"DD",X"36",X"0D",X"05",
		X"C9",X"DD",X"35",X"0A",X"DD",X"7E",X"0A",X"FE",X"50",X"D0",X"21",X"4D",X"E0",X"34",X"DD",X"36",
		X"00",X"04",X"C9",X"CD",X"DB",X"20",X"22",X"D6",X"E0",X"7C",X"D6",X"08",X"FE",X"F0",X"D2",X"52",
		X"08",X"2A",X"D8",X"E0",X"23",X"CB",X"7C",X"20",X"02",X"2B",X"2B",X"22",X"D8",X"E0",X"2A",X"DA",
		X"E0",X"ED",X"5B",X"DC",X"E0",X"19",X"4C",X"22",X"DA",X"E0",X"21",X"24",X"00",X"19",X"22",X"DC",
		X"E0",X"CB",X"14",X"38",X"1F",X"C6",X"0B",X"CD",X"38",X"15",X"D6",X"08",X"B9",X"30",X"15",X"ED",
		X"5B",X"DC",X"E0",X"21",X"00",X"00",X"ED",X"52",X"CB",X"3A",X"CB",X"1B",X"CB",X"3A",X"CB",X"1B",
		X"19",X"22",X"DC",X"E0",X"CD",X"B8",X"08",X"C3",X"EF",X"20",X"3A",X"49",X"E0",X"87",X"21",X"28",
		X"30",X"85",X"6F",X"5E",X"23",X"66",X"2E",X"00",X"22",X"0E",X"E3",X"AF",X"CB",X"13",X"17",X"57",
		X"ED",X"53",X"1C",X"E3",X"ED",X"5B",X"02",X"E3",X"AF",X"ED",X"52",X"4F",X"7C",X"30",X"03",X"ED",
		X"44",X"0C",X"FE",X"18",X"38",X"02",X"3E",X"18",X"21",X"30",X"30",X"85",X"6F",X"5E",X"16",X"00",
		X"2A",X"04",X"E3",X"7C",X"A7",X"F2",X"D4",X"14",X"0D",X"20",X"11",X"2F",X"67",X"7D",X"2F",X"6F",
		X"23",X"EB",X"18",X"03",X"0D",X"28",X"57",X"A7",X"ED",X"52",X"30",X"52",X"11",X"02",X"00",X"3A",
		X"4E",X"E0",X"1F",X"2A",X"04",X"E3",X"ED",X"5A",X"22",X"04",X"E3",X"ED",X"5B",X"02",X"E3",X"19",
		X"22",X"02",X"E3",X"54",X"21",X"DC",X"E1",X"7E",X"3D",X"C0",X"3A",X"0B",X"E5",X"87",X"87",X"87",
		X"C6",X"08",X"82",X"D0",X"36",X"00",X"21",X"0E",X"E5",X"34",X"7E",X"06",X"09",X"FE",X"19",X"28",
		X"0F",X"38",X"01",X"3D",X"D6",X"05",X"CA",X"C0",X"27",X"10",X"F9",X"FE",X"06",X"CA",X"C0",X"27",
		X"3E",X"10",X"CD",X"75",X"0D",X"AF",X"0E",X"01",X"CD",X"C2",X"02",X"C3",X"12",X"0D",X"11",X"FD",
		X"FF",X"18",X"AC",X"3A",X"03",X"E3",X"C6",X"20",X"47",X"3A",X"E2",X"E1",X"80",X"C6",X"06",X"CB",
		X"3F",X"CB",X"3F",X"6F",X"26",X"E2",X"7E",X"C9",X"2A",X"4A",X"E0",X"7C",X"AD",X"A5",X"07",X"D0",
		X"4F",X"3A",X"20",X"E3",X"A7",X"20",X"05",X"3E",X"0A",X"32",X"20",X"E3",X"21",X"30",X"E3",X"06",
		X"04",X"11",X"10",X"00",X"7E",X"A7",X"28",X"05",X"19",X"10",X"F9",X"79",X"C9",X"36",X"0E",X"3E",
		X"12",X"CD",X"75",X"0D",X"79",X"C9",X"3A",X"03",X"E3",X"4F",X"C6",X"04",X"CD",X"38",X"15",X"D6",
		X"09",X"CD",X"C9",X"15",X"7A",X"EE",X"03",X"57",X"3E",X"09",X"CD",X"92",X"15",X"2C",X"14",X"14",
		X"3E",X"0D",X"81",X"4F",X"2C",X"2C",X"7D",X"E6",X"3F",X"6F",X"7E",X"D6",X"09",X"CD",X"ED",X"08",
		X"47",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"FD",X"23",X"C3",X"76",X"09",X"3A",X"03",X"E3",X"4F",
		X"3A",X"07",X"E3",X"C6",X"11",X"CD",X"C9",X"15",X"7A",X"EE",X"03",X"57",X"3E",X"09",X"CD",X"C5",
		X"15",X"14",X"14",X"3E",X"0D",X"81",X"4F",X"18",X"D8",X"0C",X"CD",X"ED",X"08",X"47",X"11",X"00",
		X"05",X"3A",X"E2",X"E1",X"CB",X"67",X"20",X"01",X"14",X"FD",X"21",X"A4",X"E1",X"C3",X"76",X"09",
		X"DD",X"36",X"0A",X"0C",X"3A",X"07",X"E3",X"C6",X"0A",X"32",X"27",X"E3",X"2A",X"02",X"E3",X"11",
		X"00",X"1C",X"19",X"22",X"22",X"E3",X"DD",X"34",X"00",X"C9",X"DD",X"35",X"0A",X"28",X"19",X"2A",
		X"22",X"E3",X"11",X"5D",X"04",X"19",X"22",X"22",X"E3",X"DD",X"7E",X"0A",X"1F",X"3E",X"09",X"38",
		X"01",X"3C",X"DD",X"77",X"0D",X"C3",X"B8",X"08",X"DD",X"34",X"00",X"DD",X"36",X"0A",X"03",X"DD",
		X"36",X"0D",X"0B",X"3A",X"E2",X"E1",X"DD",X"86",X"03",X"DD",X"77",X"0F",X"C9",X"CD",X"31",X"08",
		X"DD",X"35",X"0A",X"F0",X"DD",X"7E",X"0D",X"FE",X"0D",X"CA",X"52",X"08",X"FE",X"29",X"CA",X"52",
		X"08",X"DD",X"34",X"0D",X"DD",X"36",X"0A",X"03",X"C9",X"3A",X"03",X"E3",X"C6",X"0A",X"DD",X"77",
		X"03",X"3A",X"07",X"E3",X"C6",X"02",X"DD",X"77",X"07",X"DD",X"34",X"00",X"C9",X"3A",X"00",X"E3",
		X"FE",X"06",X"30",X"2B",X"DD",X"7E",X"07",X"D6",X"03",X"FE",X"3A",X"38",X"22",X"DD",X"77",X"07",
		X"CD",X"1B",X"08",X"DD",X"7E",X"07",X"1F",X"1F",X"1F",X"7A",X"17",X"E6",X"07",X"F6",X"60",X"77",
		X"11",X"00",X"04",X"19",X"36",X"00",X"1F",X"D0",X"11",X"20",X"FC",X"19",X"36",X"00",X"C9",X"CD",
		X"1B",X"08",X"36",X"00",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"4E",X"03",X"DD",X"7E",X"0C",X"87",
		X"87",X"87",X"21",X"1C",X"31",X"85",X"6F",X"3A",X"20",X"E3",X"11",X"04",X"F8",X"D6",X"0B",X"28",
		X"06",X"3D",X"20",X"17",X"11",X"0A",X"F0",X"3A",X"23",X"E3",X"82",X"91",X"FE",X"E8",X"38",X"0B",
		X"3A",X"27",X"E3",X"DD",X"96",X"07",X"86",X"83",X"F2",X"4E",X"17",X"DD",X"7E",X"0C",X"A7",X"F8",
		X"23",X"3A",X"03",X"E3",X"91",X"86",X"23",X"46",X"23",X"B8",X"38",X"05",X"96",X"30",X"01",X"AF",
		X"80",X"23",X"BE",X"D2",X"C4",X"17",X"23",X"46",X"23",X"86",X"6F",X"24",X"3A",X"07",X"E3",X"86",
		X"DD",X"96",X"07",X"3D",X"80",X"F8",X"3A",X"04",X"D0",X"CB",X"77",X"C8",X"E1",X"3E",X"07",X"32",
		X"00",X"E3",X"3E",X"03",X"32",X"0D",X"E3",X"AF",X"32",X"0A",X"E3",X"32",X"B0",X"E3",X"32",X"72",
		X"E1",X"CD",X"52",X"08",X"06",X"03",X"3A",X"07",X"E3",X"C6",X"14",X"4F",X"3A",X"03",X"E3",X"21",
		X"D3",X"E1",X"34",X"21",X"C0",X"E3",X"FD",X"21",X"DF",X"30",X"36",X"1C",X"23",X"23",X"23",X"77",
		X"C6",X"10",X"CD",X"F8",X"17",X"71",X"CD",X"F8",X"17",X"23",X"23",X"FD",X"5E",X"00",X"73",X"FD",
		X"23",X"23",X"23",X"23",X"10",X"E4",X"CD",X"A1",X"08",X"3E",X"1F",X"C3",X"75",X"0D",X"3A",X"E2",
		X"E1",X"DD",X"86",X"03",X"32",X"2F",X"E3",X"3E",X"0D",X"32",X"20",X"E3",X"3E",X"26",X"32",X"2D",
		X"E3",X"3E",X"03",X"32",X"2A",X"E3",X"3E",X"01",X"CD",X"75",X"0D",X"11",X"07",X"00",X"19",X"7E",
		X"E6",X"0F",X"0E",X"01",X"FE",X"0E",X"30",X"07",X"CD",X"C2",X"02",X"E1",X"C3",X"52",X"08",X"20",
		X"13",X"CD",X"F0",X"17",X"C6",X"05",X"DD",X"77",X"08",X"CD",X"C2",X"02",X"DD",X"34",X"00",X"DD",
		X"36",X"0A",X"00",X"C9",X"CD",X"56",X"08",X"CD",X"F0",X"17",X"21",X"10",X"FB",X"C6",X"06",X"DD",
		X"77",X"08",X"E5",X"CD",X"C2",X"02",X"E1",X"DD",X"7E",X"07",X"84",X"DD",X"77",X"07",X"DD",X"7E",
		X"03",X"85",X"DD",X"77",X"03",X"DD",X"36",X"0D",X"54",X"DD",X"36",X"00",X"21",X"DD",X"36",X"0A",
		X"3B",X"C3",X"56",X"08",X"47",X"DD",X"7E",X"0C",X"C6",X"80",X"4F",X"FE",X"8B",X"28",X"1B",X"FE",
		X"8E",X"28",X"17",X"78",X"96",X"FE",X"04",X"D0",X"DD",X"71",X"0C",X"23",X"23",X"23",X"7E",X"1F",
		X"1F",X"1F",X"1F",X"E6",X"0F",X"0E",X"01",X"C3",X"C2",X"02",X"78",X"FE",X"FC",X"30",X"E9",X"C9",
		X"ED",X"5F",X"E6",X"03",X"C0",X"3E",X"02",X"C9",X"23",X"FD",X"5E",X"00",X"73",X"23",X"FD",X"5E",
		X"01",X"73",X"23",X"23",X"FD",X"23",X"FD",X"23",X"C9",X"3A",X"00",X"E3",X"FE",X"06",X"D0",X"FE",
		X"01",X"26",X"00",X"28",X"76",X"2A",X"1C",X"E3",X"ED",X"5B",X"1A",X"E3",X"7A",X"A7",X"FA",X"23",
		X"18",X"ED",X"52",X"21",X"03",X"00",X"30",X"03",X"21",X"FE",X"FF",X"3A",X"4E",X"E0",X"1F",X"38",
		X"01",X"1D",X"19",X"22",X"1A",X"E3",X"ED",X"5B",X"04",X"E3",X"A7",X"ED",X"52",X"22",X"14",X"E3",
		X"EB",X"2A",X"E1",X"E1",X"19",X"22",X"E1",X"E1",X"3A",X"D9",X"E1",X"1F",X"30",X"3D",X"2A",X"EF",
		X"E0",X"19",X"7C",X"C6",X"06",X"FE",X"0C",X"38",X"17",X"D6",X"12",X"67",X"E5",X"21",X"3F",X"E2",
		X"11",X"42",X"E2",X"01",X"40",X"00",X"ED",X"B8",X"21",X"42",X"E2",X"0E",X"03",X"ED",X"B8",X"E1",
		X"22",X"EF",X"E0",X"ED",X"5B",X"F1",X"E0",X"19",X"3A",X"08",X"E5",X"FE",X"03",X"30",X"0C",X"3A",
		X"E2",X"E1",X"94",X"FE",X"F4",X"38",X"04",X"AF",X"32",X"D9",X"E1",X"7C",X"2F",X"21",X"3D",X"E0",
		X"86",X"32",X"C0",X"E1",X"2A",X"14",X"E3",X"54",X"5D",X"CB",X"3C",X"CB",X"1D",X"19",X"CB",X"3C",
		X"CB",X"1D",X"CB",X"3C",X"CB",X"1D",X"EB",X"2A",X"04",X"E5",X"19",X"22",X"04",X"E5",X"7C",X"2F",
		X"32",X"C1",X"E1",X"CB",X"3A",X"CB",X"1B",X"2A",X"06",X"E5",X"19",X"22",X"06",X"E5",X"7C",X"2F",
		X"32",X"C2",X"E1",X"CD",X"33",X"15",X"FE",X"C4",X"30",X"02",X"3E",X"C4",X"C6",X"28",X"30",X"01",
		X"AF",X"47",X"C6",X"94",X"32",X"C3",X"E1",X"CB",X"28",X"78",X"C6",X"72",X"32",X"C4",X"E1",X"C9",
		X"CD",X"31",X"08",X"CD",X"99",X"16",X"DD",X"35",X"0A",X"F0",X"DD",X"34",X"0A",X"DD",X"7E",X"03",
		X"FE",X"E0",X"D0",X"DD",X"7E",X"0C",X"17",X"D8",X"3A",X"C0",X"E3",X"A7",X"C0",X"FD",X"21",X"70",
		X"E3",X"11",X"10",X"00",X"06",X"05",X"FD",X"7E",X"00",X"FE",X"1D",X"20",X"0D",X"FD",X"7E",X"0C",
		X"17",X"38",X"07",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"D8",X"FD",X"19",X"10",X"E8",X"DD",X"7E",
		X"07",X"FD",X"77",X"07",X"DD",X"7E",X"0F",X"D6",X"04",X"FD",X"77",X"0F",X"FD",X"36",X"00",X"11",
		X"FD",X"36",X"0D",X"22",X"FD",X"36",X"0C",X"0C",X"DD",X"36",X"0A",X"43",X"C9",X"3A",X"00",X"E3",
		X"FE",X"06",X"D0",X"DD",X"7E",X"04",X"C6",X"DD",X"DD",X"77",X"04",X"30",X"03",X"DD",X"35",X"0F",
		X"CD",X"38",X"08",X"CD",X"99",X"16",X"C9",X"CD",X"31",X"08",X"CD",X"99",X"16",X"C9",X"CD",X"31",
		X"08",X"DD",X"7E",X"0C",X"A7",X"C0",X"DD",X"7E",X"0D",X"07",X"07",X"E6",X"1C",X"21",X"00",X"2E",
		X"85",X"6F",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"86",X"23",X"BE",X"30",X"45",X"47",X"3A",X"00",
		X"E3",X"FE",X"04",X"C8",X"3A",X"04",X"D0",X"CB",X"77",X"C8",X"78",X"46",X"0E",X"02",X"CB",X"38",
		X"50",X"CB",X"38",X"BA",X"38",X"04",X"78",X"82",X"47",X"0D",X"DD",X"7E",X"03",X"80",X"D6",X"1C",
		X"32",X"03",X"E3",X"79",X"32",X"0D",X"E3",X"3D",X"3D",X"32",X"05",X"E3",X"3E",X"80",X"32",X"04",
		X"E3",X"23",X"7E",X"32",X"0A",X"E3",X"21",X"00",X"02",X"22",X"08",X"E3",X"3E",X"06",X"32",X"00",
		X"E3",X"C9",X"96",X"FE",X"04",X"D0",X"DD",X"34",X"0C",X"23",X"23",X"7E",X"0E",X"01",X"C3",X"C2",
		X"02",X"DD",X"35",X"0A",X"F2",X"0D",X"1A",X"DD",X"7E",X"0E",X"47",X"3C",X"0E",X"07",X"FE",X"06",
		X"38",X"0B",X"3A",X"4E",X"E0",X"E6",X"30",X"20",X"02",X"3E",X"30",X"4F",X"AF",X"DD",X"77",X"0E",
		X"DD",X"71",X"0A",X"78",X"FE",X"04",X"38",X"04",X"EE",X"07",X"3D",X"47",X"C6",X"06",X"DD",X"46",
		X"0C",X"04",X"FA",X"08",X"1A",X"DD",X"77",X"0C",X"C6",X"45",X"DD",X"77",X"0D",X"3A",X"20",X"E3",
		X"FE",X"0F",X"38",X"0E",X"C0",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"C6",X"10",X"FE",X"30",X"DA",
		X"FD",X"16",X"CD",X"38",X"08",X"DD",X"7E",X"0C",X"FE",X"06",X"C8",X"CD",X"99",X"16",X"C9",X"CD",
		X"31",X"08",X"DD",X"35",X"0A",X"F0",X"DD",X"7E",X"0D",X"FE",X"4A",X"C8",X"DD",X"35",X"0D",X"DD",
		X"36",X"0A",X"07",X"C9",X"3A",X"00",X"E3",X"FE",X"06",X"D0",X"DD",X"35",X"0E",X"F2",X"66",X"1A",
		X"DD",X"36",X"0E",X"06",X"DD",X"7E",X"0D",X"3D",X"01",X"03",X"00",X"21",X"8E",X"1A",X"ED",X"B1",
		X"20",X"01",X"7E",X"DD",X"77",X"0D",X"DD",X"7E",X"04",X"C6",X"C0",X"DD",X"77",X"04",X"30",X"03",
		X"DD",X"35",X"0F",X"CD",X"38",X"08",X"DD",X"7E",X"0C",X"D6",X"04",X"CB",X"27",X"C6",X"0C",X"4F",
		X"DD",X"7E",X"03",X"CD",X"38",X"15",X"91",X"DD",X"77",X"07",X"CD",X"99",X"16",X"C9",X"11",X"15",
		X"1A",X"20",X"DD",X"36",X"0B",X"01",X"3A",X"00",X"E3",X"FE",X"06",X"D0",X"2A",X"72",X"E3",X"7C",
		X"FE",X"08",X"28",X"09",X"11",X"70",X"00",X"19",X"22",X"72",X"E3",X"18",X"2C",X"DD",X"36",X"0A",
		X"00",X"DD",X"34",X"00",X"DD",X"36",X"0E",X"80",X"C9",X"3A",X"4E",X"E0",X"1F",X"D8",X"3A",X"00",
		X"E3",X"FE",X"06",X"D0",X"3A",X"4E",X"E0",X"47",X"E6",X"03",X"20",X"0D",X"DD",X"34",X"03",X"CB",
		X"68",X"28",X"06",X"DD",X"35",X"03",X"DD",X"35",X"03",X"3A",X"4E",X"E0",X"E6",X"07",X"20",X"0D",
		X"DD",X"7E",X"03",X"C6",X"18",X"CD",X"38",X"15",X"D6",X"10",X"DD",X"77",X"07",X"C3",X"B8",X"08",
		X"DD",X"35",X"0E",X"20",X"CF",X"DD",X"36",X"0A",X"58",X"DD",X"34",X"00",X"DD",X"36",X"0D",X"52",
		X"C9",X"DD",X"35",X"0A",X"28",X"15",X"2A",X"72",X"E3",X"11",X"80",X"01",X"19",X"22",X"72",X"E3",
		X"7C",X"FE",X"F0",X"D2",X"52",X"08",X"CD",X"99",X"16",X"18",X"BE",X"DD",X"34",X"00",X"DD",X"36",
		X"0A",X"6E",X"DD",X"36",X"0D",X"23",X"C9",X"CD",X"99",X"16",X"DD",X"35",X"0A",X"20",X"95",X"DD",
		X"35",X"00",X"DD",X"35",X"0B",X"DD",X"36",X"0D",X"52",X"C9",X"21",X"EE",X"E0",X"3A",X"4E",X"E0",
		X"96",X"F8",X"01",X"00",X"10",X"ED",X"5F",X"E6",X"F0",X"26",X"E4",X"51",X"59",X"6F",X"7E",X"D6",
		X"1E",X"FE",X"0A",X"30",X"0A",X"CB",X"4F",X"20",X"06",X"FE",X"04",X"38",X"63",X"0C",X"5D",X"7D",
		X"C6",X"10",X"10",X"E9",X"ED",X"53",X"D4",X"E1",X"0D",X"F8",X"3A",X"10",X"E5",X"E6",X"03",X"FE",
		X"01",X"89",X"4F",X"FE",X"09",X"DA",X"7A",X"1B",X"0E",X"08",X"21",X"FF",X"2F",X"09",X"4E",X"06",
		X"05",X"21",X"70",X"E3",X"11",X"00",X"00",X"7E",X"A7",X"28",X"39",X"D6",X"2F",X"20",X"01",X"14",
		X"7D",X"C6",X"10",X"6F",X"10",X"F1",X"7A",X"B9",X"D0",X"1C",X"1D",X"C8",X"ED",X"5F",X"E6",X"0F",
		X"C6",X"19",X"21",X"4E",X"E0",X"86",X"32",X"EE",X"E0",X"16",X"00",X"DD",X"21",X"00",X"E3",X"DD",
		X"19",X"21",X"D4",X"E1",X"5E",X"FD",X"21",X"00",X"E4",X"FD",X"19",X"0E",X"3B",X"C3",X"64",X"10",
		X"55",X"14",X"18",X"9B",X"5D",X"18",X"C9",X"3A",X"4E",X"E0",X"21",X"52",X"E0",X"AE",X"E6",X"1F",
		X"C0",X"ED",X"5F",X"77",X"21",X"C6",X"E1",X"06",X"03",X"7E",X"A7",X"20",X"04",X"23",X"10",X"F9",
		X"C9",X"DD",X"21",X"00",X"E4",X"04",X"78",X"48",X"06",X"10",X"FE",X"04",X"28",X"0F",X"3A",X"D6",
		X"E1",X"3D",X"FA",X"FD",X"1B",X"0D",X"0D",X"DD",X"21",X"70",X"E3",X"06",X"05",X"11",X"10",X"00",
		X"DD",X"7E",X"00",X"A7",X"28",X"05",X"DD",X"19",X"10",X"F6",X"C9",X"35",X"79",X"FE",X"02",X"30",
		X"43",X"ED",X"5F",X"E6",X"1F",X"C6",X"20",X"DD",X"77",X"0F",X"21",X"D6",X"E1",X"35",X"ED",X"5F",
		X"E6",X"1E",X"5F",X"16",X"00",X"FE",X"0E",X"3E",X"82",X"38",X"04",X"ED",X"5F",X"E6",X"80",X"DD",
		X"77",X"0C",X"21",X"08",X"30",X"19",X"7E",X"DD",X"77",X"07",X"23",X"7E",X"DD",X"77",X"03",X"06",
		X"00",X"21",X"59",X"1C",X"09",X"09",X"7E",X"DD",X"77",X"0D",X"DD",X"36",X"0E",X"00",X"23",X"7E",
		X"DD",X"77",X"00",X"C9",X"CD",X"0A",X"08",X"18",X"C5",X"2B",X"26",X"2A",X"26",X"2B",X"22",X"2A",
		X"22",X"31",X"1E",X"DD",X"7E",X"0D",X"FE",X"2B",X"D8",X"DD",X"CB",X"0E",X"7E",X"20",X"18",X"DD",
		X"35",X"0E",X"F0",X"DD",X"34",X"0D",X"FE",X"2F",X"28",X"1C",X"FE",X"34",X"20",X"04",X"DD",X"36",
		X"0D",X"31",X"DD",X"36",X"0E",X"08",X"C9",X"DD",X"34",X"0E",X"F8",X"DD",X"35",X"0D",X"FE",X"2C",
		X"28",X"F0",X"FE",X"32",X"28",X"EC",X"DD",X"36",X"0E",X"F8",X"C9",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"CB",X"3C",X"CB",X"1D",X"DD",X"CB",X"0C",X"46",X"28",X"07",X"EB",X"21",X"00",X"00",X"A7",
		X"ED",X"52",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",X"34",X"00",X"C9",X"0E",X"3D",X"DD",X"7E",
		X"09",X"A7",X"20",X"13",X"0E",X"3B",X"DD",X"46",X"05",X"CB",X"10",X"30",X"02",X"0E",X"50",X"DD",
		X"7E",X"08",X"FE",X"60",X"38",X"01",X"0C",X"DD",X"71",X"0D",X"CD",X"FB",X"20",X"7C",X"FE",X"06",
		X"DA",X"52",X"08",X"01",X"05",X"00",X"22",X"D6",X"E0",X"7C",X"2A",X"DC",X"E0",X"09",X"22",X"DC",
		X"E0",X"ED",X"5B",X"DA",X"E0",X"19",X"22",X"DA",X"E0",X"54",X"CD",X"38",X"15",X"D6",X"08",X"BA",
		X"CD",X"EF",X"20",X"30",X"35",X"DD",X"77",X"07",X"DD",X"34",X"00",X"DD",X"36",X"0B",X"00",X"DD",
		X"7E",X"00",X"FE",X"2A",X"3E",X"03",X"20",X"05",X"DD",X"36",X"00",X"30",X"3D",X"CD",X"75",X"0D",
		X"C3",X"56",X"08",X"CD",X"DB",X"20",X"ED",X"5B",X"14",X"E3",X"CB",X"2A",X"CB",X"1B",X"ED",X"52",
		X"11",X"8E",X"00",X"ED",X"52",X"01",X"10",X"00",X"18",X"AC",X"3A",X"00",X"E3",X"FE",X"06",X"D2",
		X"B8",X"08",X"21",X"05",X"06",X"DD",X"7E",X"00",X"FE",X"2A",X"30",X"03",X"21",X"0B",X"02",X"FD",
		X"21",X"30",X"E3",X"11",X"10",X"00",X"06",X"04",X"FD",X"7E",X"00",X"FE",X"0F",X"20",X"14",X"FD",
		X"7E",X"07",X"DD",X"96",X"07",X"FE",X"0A",X"30",X"0A",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"94",
		X"BD",X"38",X"2B",X"FD",X"19",X"10",X"E1",X"3A",X"07",X"E3",X"DD",X"96",X"07",X"FE",X"F0",X"DA",
		X"B8",X"08",X"57",X"3A",X"03",X"E3",X"DD",X"96",X"03",X"D6",X"04",X"FE",X"EA",X"DA",X"B8",X"08",
		X"3A",X"04",X"D0",X"CB",X"77",X"CA",X"B8",X"08",X"CD",X"52",X"08",X"C3",X"FD",X"16",X"FD",X"34",
		X"00",X"DD",X"7E",X"0D",X"FE",X"37",X"38",X"11",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"00",X"2D",
		X"DD",X"36",X"0A",X"0A",X"DD",X"36",X"0D",X"4F",X"C9",X"21",X"C9",X"E1",X"01",X"01",X"05",X"FE",
		X"31",X"30",X"07",X"23",X"05",X"FE",X"2A",X"28",X"01",X"23",X"3E",X"11",X"CD",X"75",X"0D",X"35",
		X"20",X"08",X"23",X"23",X"23",X"7E",X"FE",X"03",X"30",X"11",X"DD",X"36",X"00",X"20",X"DD",X"36",
		X"0A",X"06",X"DD",X"36",X"0D",X"37",X"78",X"CD",X"C2",X"02",X"C9",X"21",X"00",X"FC",X"D6",X"02",
		X"C3",X"9D",X"17",X"DD",X"36",X"0D",X"3E",X"CD",X"23",X"16",X"D6",X"03",X"E6",X"F8",X"C6",X"06",
		X"DD",X"77",X"0F",X"21",X"D1",X"E1",X"7E",X"A7",X"28",X"13",X"23",X"36",X"01",X"23",X"7E",X"A7",
		X"C8",X"C3",X"52",X"08",X"DD",X"36",X"0D",X"43",X"CD",X"23",X"16",X"18",X"E6",X"34",X"DD",X"34",
		X"00",X"DD",X"36",X"0A",X"04",X"CD",X"31",X"08",X"C9",X"21",X"D2",X"E1",X"7E",X"23",X"B6",X"A7",
		X"C2",X"52",X"08",X"DD",X"7E",X"03",X"FE",X"F8",X"D2",X"52",X"08",X"DD",X"35",X"0A",X"20",X"E5",
		X"DD",X"7E",X"0D",X"FE",X"49",X"CA",X"52",X"08",X"DD",X"34",X"0D",X"DD",X"36",X"0A",X"05",X"18",
		X"D4",X"3A",X"D3",X"E1",X"A7",X"C2",X"52",X"08",X"DD",X"35",X"0A",X"20",X"C8",X"DD",X"7E",X"0D",
		X"FE",X"42",X"30",X"1F",X"DD",X"34",X"0D",X"FE",X"3F",X"20",X"12",X"DD",X"7E",X"0F",X"1F",X"1F",
		X"1F",X"E6",X"1F",X"5F",X"16",X"83",X"0E",X"09",X"3E",X"01",X"CD",X"C2",X"02",X"DD",X"36",X"0A",
		X"02",X"18",X"A2",X"DD",X"7E",X"07",X"C6",X"08",X"DD",X"77",X"07",X"CD",X"56",X"08",X"DD",X"36",
		X"0C",X"00",X"DD",X"36",X"0D",X"81",X"DD",X"36",X"00",X"13",X"C9",X"DD",X"35",X"0A",X"CA",X"52",
		X"08",X"C3",X"B8",X"08",X"DD",X"35",X"0F",X"CA",X"4D",X"20",X"DD",X"34",X"00",X"DD",X"7E",X"0C",
		X"CB",X"27",X"28",X"3D",X"3F",X"1F",X"E6",X"80",X"DD",X"77",X"0C",X"4F",X"ED",X"5F",X"E6",X"3F",
		X"5F",X"16",X"00",X"21",X"26",X"01",X"19",X"0C",X"F2",X"D2",X"1E",X"EB",X"A7",X"21",X"00",X"00",
		X"ED",X"52",X"DD",X"74",X"05",X"DD",X"75",X"04",X"EE",X"3F",X"D6",X"20",X"87",X"DD",X"77",X"08",
		X"3E",X"00",X"DE",X"00",X"DD",X"77",X"09",X"ED",X"5F",X"E6",X"7F",X"C6",X"20",X"DD",X"77",X"0A",
		X"C9",X"06",X"01",X"DD",X"7E",X"07",X"FE",X"44",X"38",X"0C",X"06",X"03",X"FE",X"58",X"30",X"06",
		X"ED",X"5F",X"E6",X"02",X"3C",X"47",X"78",X"DD",X"86",X"0C",X"DD",X"77",X"0C",X"ED",X"5F",X"E6",
		X"0F",X"C6",X"24",X"DD",X"77",X"0B",X"21",X"66",X"01",X"DD",X"75",X"04",X"DD",X"74",X"05",X"DD",
		X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"C9",X"CD",X"63",X"1C",X"CD",X"DB",X"20",X"DD",X"7E",
		X"0C",X"CB",X"27",X"20",X"52",X"DD",X"35",X"0A",X"28",X"49",X"2A",X"D6",X"E0",X"ED",X"5B",X"D8",
		X"E0",X"19",X"7A",X"ED",X"5B",X"04",X"E3",X"ED",X"52",X"22",X"D6",X"E0",X"17",X"38",X"2F",X"DD",
		X"7E",X"0D",X"06",X"A0",X"D6",X"2A",X"28",X"08",X"06",X"80",X"D6",X"07",X"38",X"02",X"06",X"D0",
		X"7C",X"B8",X"30",X"1F",X"2A",X"DA",X"E0",X"ED",X"5B",X"DC",X"E0",X"19",X"22",X"DA",X"E0",X"7C",
		X"FE",X"38",X"38",X"0F",X"FE",X"70",X"30",X"0B",X"CD",X"EF",X"20",X"C3",X"4C",X"1D",X"7C",X"FE",
		X"16",X"30",X"E1",X"DD",X"35",X"00",X"C9",X"2A",X"D8",X"E0",X"DD",X"5E",X"0B",X"16",X"00",X"A7",
		X"ED",X"52",X"22",X"D8",X"E0",X"30",X"16",X"DD",X"7E",X"03",X"D6",X"30",X"FE",X"40",X"3E",X"00",
		X"30",X"04",X"ED",X"5F",X"E6",X"80",X"DD",X"86",X"0C",X"3C",X"DD",X"77",X"0C",X"EB",X"2A",X"D6",
		X"E0",X"ED",X"52",X"DD",X"7E",X"0C",X"07",X"38",X"02",X"19",X"19",X"ED",X"5B",X"04",X"E3",X"ED",
		X"52",X"22",X"D6",X"E0",X"2A",X"DC",X"E0",X"DD",X"5E",X"0B",X"16",X"00",X"0F",X"3D",X"0F",X"30",
		X"1A",X"A7",X"ED",X"52",X"38",X"AD",X"22",X"DC",X"E0",X"EB",X"2A",X"DA",X"E0",X"A7",X"ED",X"52",
		X"0F",X"38",X"02",X"19",X"19",X"22",X"DA",X"E0",X"C3",X"78",X"1F",X"19",X"18",X"E8",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"34",X"00",X"DD",X"7E",X"0C",X"E6",X"7F",X"C8",X"CD",X"28",X"1F",X"DD",X"7E",X"00",X"FE",
		X"25",X"CA",X"83",X"1F",X"FE",X"24",X"CA",X"AA",X"1E",X"C9",X"CD",X"63",X"1C",X"CD",X"DB",X"20",
		X"22",X"D6",X"E0",X"7C",X"D6",X"08",X"FE",X"F0",X"D2",X"52",X"08",X"ED",X"5B",X"DC",X"E0",X"2A",
		X"DA",X"E0",X"19",X"22",X"DA",X"E0",X"7C",X"FE",X"30",X"DA",X"52",X"08",X"7A",X"A7",X"FA",X"78",
		X"1F",X"21",X"00",X"00",X"A7",X"ED",X"52",X"22",X"DC",X"E0",X"C3",X"78",X"1F",X"3A",X"03",X"E3",
		X"16",X"00",X"C6",X"10",X"DD",X"96",X"03",X"30",X"03",X"ED",X"44",X"15",X"1F",X"1F",X"1F",X"E6",
		X"1E",X"4F",X"06",X"00",X"21",X"24",X"2D",X"09",X"FE",X"12",X"38",X"01",X"04",X"7E",X"CB",X"7A",
		X"28",X"06",X"2F",X"5F",X"78",X"2F",X"47",X"7B",X"DD",X"77",X"04",X"DD",X"70",X"05",X"23",X"5E",
		X"16",X"00",X"79",X"FE",X"0A",X"30",X"01",X"14",X"DD",X"72",X"09",X"DD",X"73",X"08",X"DD",X"36",
		X"00",X"29",X"2A",X"1A",X"E3",X"DD",X"75",X"0B",X"DD",X"74",X"0F",X"C9",X"CD",X"63",X"1C",X"CD",
		X"FB",X"20",X"22",X"D6",X"E0",X"7C",X"2A",X"DC",X"E0",X"C3",X"F1",X"1C",X"DD",X"35",X"0A",X"C2",
		X"B8",X"08",X"DD",X"36",X"0A",X"06",X"DD",X"7E",X"0D",X"FE",X"39",X"D2",X"52",X"08",X"DD",X"34",
		X"0D",X"C3",X"B8",X"08",X"DD",X"35",X"0A",X"C2",X"B8",X"08",X"DD",X"7E",X"07",X"FE",X"80",X"D2",
		X"52",X"08",X"06",X"80",X"DD",X"36",X"00",X"00",X"C3",X"69",X"08",X"DD",X"E5",X"E1",X"11",X"D4",
		X"E0",X"01",X"0A",X"00",X"ED",X"B0",X"ED",X"5B",X"D6",X"E0",X"2A",X"D8",X"E0",X"19",X"C9",X"DD",
		X"E5",X"D1",X"21",X"D4",X"E0",X"01",X"0A",X"00",X"ED",X"B0",X"C9",X"CD",X"DB",X"20",X"EB",X"DD",
		X"6E",X"0B",X"DD",X"66",X"0F",X"ED",X"4B",X"1A",X"E3",X"ED",X"42",X"19",X"C9",X"21",X"51",X"E0",
		X"3A",X"00",X"E3",X"3D",X"28",X"11",X"7E",X"A7",X"F0",X"21",X"11",X"E5",X"3E",X"01",X"86",X"27",
		X"77",X"23",X"7E",X"CE",X"00",X"27",X"77",X"3E",X"37",X"32",X"51",X"E0",X"11",X"90",X"80",X"FD",
		X"21",X"90",X"84",X"0E",X"02",X"CD",X"E7",X"03",X"3A",X"12",X"E5",X"CD",X"BD",X"03",X"3A",X"11",
		X"E5",X"C3",X"AE",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"01",X"03",X"34",X"07",X"49",X"08",X"63",X"0F",X"73",X"07",X"80",X"19",X"92",X"0F",
		X"A0",X"06",X"A1",X"03",X"A2",X"2A",X"E0",X"32",X"FF",X"28",X"0F",X"0F",X"3F",X"30",X"40",X"06",
		X"41",X"03",X"42",X"2A",X"4C",X"0F",X"92",X"0F",X"9F",X"28",X"A5",X"07",X"B8",X"0F",X"CD",X"0F",
		X"E0",X"06",X"E1",X"03",X"00",X"19",X"01",X"08",X"14",X"07",X"20",X"33",X"4F",X"0F",X"7F",X"30",
		X"80",X"06",X"81",X"03",X"82",X"22",X"9C",X"1C",X"B6",X"1C",X"C0",X"2A",X"D9",X"1C",X"DF",X"20",
		X"03",X"0F",X"08",X"28",X"16",X"07",X"20",X"06",X"21",X"03",X"3C",X"22",X"52",X"1C",X"60",X"32",
		X"6E",X"1C",X"7F",X"20",X"A6",X"08",X"B7",X"0F",X"BF",X"30",X"C0",X"06",X"C1",X"03",X"C4",X"08",
		X"D3",X"0A",X"E6",X"0E",X"F6",X"0F",X"0C",X"10",X"1C",X"0F",X"2D",X"0E",X"39",X"07",X"4A",X"0F",
		X"5B",X"0F",X"60",X"06",X"61",X"03",X"6E",X"19",X"6F",X"09",X"82",X"0F",X"8F",X"09",X"A0",X"2B",
		X"A2",X"0F",X"B1",X"0F",X"FF",X"28",X"00",X"06",X"01",X"03",X"02",X"22",X"14",X"1C",X"28",X"1C",
		X"40",X"2A",X"54",X"1C",X"5F",X"20",X"9F",X"28",X"A0",X"06",X"A1",X"03",X"A2",X"23",X"A6",X"1C",
		X"D3",X"1C",X"E9",X"0F",X"F7",X"0A",X"FF",X"20",X"07",X"10",X"17",X"0E",X"29",X"10",X"35",X"0A",
		X"40",X"06",X"41",X"02",X"42",X"1A",X"60",X"03",X"6F",X"12",X"78",X"12",X"88",X"12",X"92",X"12",
		X"A3",X"12",X"A4",X"12",X"B1",X"12",X"C2",X"12",X"CD",X"12",X"CE",X"12",X"D9",X"12",X"E0",X"06",
		X"E1",X"03",X"EB",X"12",X"FA",X"12",X"06",X"12",X"07",X"12",X"14",X"12",X"23",X"12",X"2C",X"12",
		X"37",X"12",X"42",X"12",X"56",X"12",X"57",X"12",X"65",X"12",X"6E",X"12",X"7A",X"12",X"80",X"06",
		X"81",X"03",X"85",X"12",X"86",X"12",X"91",X"12",X"92",X"12",X"A3",X"12",X"A4",X"12",X"AE",X"12",
		X"B8",X"12",X"B9",X"12",X"CA",X"12",X"CB",X"12",X"D7",X"12",X"E3",X"12",X"F3",X"12",X"00",X"19",
		X"20",X"06",X"21",X"03",X"22",X"2C",X"60",X"33",X"9F",X"28",X"BF",X"30",X"C0",X"06",X"C1",X"03",
		X"C2",X"24",X"D5",X"1C",X"EA",X"1C",X"00",X"33",X"05",X"1C",X"18",X"1C",X"31",X"1C",X"3F",X"20",
		X"48",X"30",X"60",X"06",X"61",X"03",X"7B",X"24",X"87",X"1C",X"99",X"1C",X"A0",X"2B",X"AE",X"1C",
		X"C5",X"1C",X"D7",X"1C",X"DF",X"20",X"E0",X"28",X"00",X"06",X"01",X"04",X"13",X"14",X"1E",X"16",
		X"2D",X"16",X"2F",X"16",X"3A",X"15",X"4C",X"16",X"4E",X"16",X"58",X"16",X"66",X"16",X"68",X"16",
		X"72",X"02",X"73",X"14",X"7E",X"16",X"80",X"19",X"A0",X"86",X"A1",X"03",X"A2",X"34",X"C7",X"0F",
		X"EC",X"10",X"0F",X"0A",X"1F",X"30",X"2A",X"10",X"40",X"86",X"41",X"02",X"42",X"19",X"60",X"32",
		X"61",X"05",X"80",X"2A",X"BF",X"30",X"C0",X"02",X"DF",X"28",X"E0",X"06",X"E1",X"03",X"E2",X"2B",
		X"00",X"23",X"01",X"03",X"2A",X"1C",X"3F",X"28",X"45",X"1C",X"57",X"1C",X"6C",X"1C",X"6D",X"20",
		X"80",X"06",X"81",X"02",X"A0",X"03",X"A8",X"10",X"B4",X"0A",X"C5",X"07",X"DC",X"0F",X"E3",X"09",
		X"F2",X"07",X"0A",X"10",X"0D",X"09",X"1C",X"08",X"20",X"06",X"21",X"03",X"2C",X"0F",X"2F",X"0F",
		X"32",X"0A",X"45",X"13",X"54",X"13",X"66",X"13",X"77",X"0A",X"8A",X"13",X"98",X"13",X"A7",X"13",
		X"B4",X"13",X"C0",X"06",X"C1",X"03",X"C5",X"09",X"D4",X"0A",X"E0",X"02",X"E7",X"0A",X"F5",X"09",
		X"00",X"04",X"1C",X"16",X"2A",X"15",X"2C",X"15",X"35",X"16",X"3D",X"14",X"40",X"02",X"48",X"14",
		X"4A",X"14",X"60",X"86",X"61",X"02",X"62",X"19",X"80",X"03",X"81",X"2C",X"A0",X"33",X"DF",X"28",
		X"FF",X"30",X"00",X"86",X"01",X"03",X"02",X"2C",X"40",X"23",X"57",X"1C",X"5F",X"28",X"6C",X"1C",
		X"83",X"1C",X"9A",X"1C",X"A0",X"86",X"A1",X"03",X"A2",X"23",X"AE",X"1C",X"C5",X"1C",X"D5",X"1C",
		X"E0",X"33",X"E8",X"1C",X"F5",X"0F",X"FF",X"20",X"0A",X"09",X"1C",X"0A",X"28",X"30",X"32",X"10",
		X"40",X"06",X"42",X"02",X"5B",X"2B",X"60",X"03",X"80",X"33",X"9F",X"28",X"D0",X"30",X"E0",X"06",
		X"E1",X"03",X"E2",X"1B",X"20",X"17",X"60",X"18",X"80",X"06",X"81",X"03",X"C6",X"13",X"D2",X"0F",
		X"DD",X"0F",X"EE",X"0E",X"FC",X"0A",X"01",X"13",X"0D",X"09",X"20",X"06",X"21",X"03",X"22",X"13",
		X"2B",X"13",X"39",X"13",X"49",X"13",X"4C",X"0A",X"5C",X"0F",X"6A",X"0F",X"79",X"13",X"84",X"13",
		X"86",X"0A",X"95",X"0F",X"A4",X"13",X"B3",X"13",X"B5",X"09",X"C0",X"06",X"C1",X"02",X"C2",X"19",
		X"E0",X"03",X"E1",X"2C",X"EA",X"07",X"F9",X"09",X"07",X"0A",X"19",X"0F",X"2A",X"0F",X"39",X"09",
		X"48",X"28",X"54",X"0F",X"60",X"06",X"61",X"03",X"7B",X"23",X"84",X"1C",X"92",X"1C",X"A0",X"23",
		X"A3",X"1C",X"B3",X"1C",X"C3",X"1C",X"DC",X"1C",X"EF",X"1C",X"FF",X"20",X"00",X"06",X"01",X"03",
		X"07",X"10",X"0A",X"0A",X"1A",X"0F",X"2C",X"09",X"32",X"0F",X"41",X"07",X"4F",X"08",X"5C",X"0F",
		X"63",X"09",X"70",X"07",X"7D",X"0E",X"80",X"19",X"A0",X"06",X"A1",X"03",X"A2",X"24",X"AF",X"1C",
		X"BC",X"1C",X"C0",X"2C",X"CA",X"1C",X"D9",X"1C",X"E8",X"1C",X"F6",X"1C",X"FF",X"28",X"05",X"0A",
		X"10",X"1C",X"11",X"20",X"25",X"0C",X"32",X"0F",X"35",X"0C",X"40",X"06",X"41",X"03",X"42",X"19",
		X"60",X"33",X"80",X"2B",X"83",X"0A",X"92",X"07",X"BF",X"30",X"C6",X"0F",X"C9",X"0A",X"D9",X"09",
		X"DF",X"28",X"E0",X"06",X"E1",X"03",X"E2",X"24",X"EA",X"1C",X"04",X"0A",X"14",X"0F",X"1C",X"1C",
		X"24",X"20",X"34",X"09",X"45",X"0F",X"49",X"0F",X"4B",X"0C",X"58",X"0C",X"67",X"0C",X"75",X"0C",
		X"7A",X"0F",X"80",X"06",X"81",X"02",X"90",X"04",X"AD",X"16",X"B7",X"15",X"BE",X"14",X"C5",X"16",
		X"C7",X"16",X"D4",X"14",X"DB",X"15",X"E6",X"14",X"E8",X"14",X"E9",X"16",X"F0",X"14",X"F1",X"16",
		X"F2",X"14",X"02",X"15",X"04",X"15",X"0E",X"16",X"0F",X"02",X"10",X"14",X"13",X"16",X"17",X"14",
		X"19",X"14",X"20",X"86",X"21",X"03",X"22",X"19",X"40",X"2C",X"41",X"33",X"42",X"03",X"BE",X"28",
		X"BF",X"30",X"C0",X"86",X"C1",X"03",X"C2",X"1A",X"E8",X"12",X"F2",X"12",X"F4",X"12",X"FD",X"12",
		X"08",X"12",X"13",X"12",X"22",X"12",X"23",X"12",X"2E",X"12",X"36",X"12",X"42",X"12",X"4E",X"12",
		X"57",X"12",X"60",X"86",X"61",X"03",X"65",X"12",X"67",X"12",X"72",X"12",X"7A",X"12",X"83",X"12",
		X"8F",X"12",X"97",X"12",X"A2",X"12",X"AB",X"12",X"B7",X"12",X"C2",X"12",X"D0",X"12",X"D8",X"12",
		X"E4",X"12",X"00",X"86",X"01",X"03",X"20",X"25",X"25",X"09",X"33",X"1C",X"40",X"2C",X"48",X"10",
		X"54",X"1C",X"65",X"0F",X"6F",X"1C",X"7F",X"20",X"80",X"02",X"88",X"28",X"A0",X"86",X"A1",X"05",
		X"BB",X"35",X"C0",X"2C",X"DF",X"02",X"FF",X"30",X"0A",X"10",X"19",X"0A",X"1F",X"28",X"20",X"03",
		X"29",X"0F",X"2C",X"0A",X"32",X"0F",X"3A",X"0F",X"40",X"06",X"41",X"02",X"47",X"0F",X"4A",X"0A",
		X"50",X"0F",X"60",X"03",X"65",X"07",X"79",X"08",X"80",X"17",X"8A",X"0A",X"A0",X"18",X"C8",X"09",
		X"E0",X"06",X"E1",X"03",X"EF",X"10",X"F4",X"0F",X"F7",X"0A",X"06",X"0F",X"11",X"10",X"14",X"09",
		X"1A",X"1A",X"3A",X"12",X"42",X"12",X"44",X"12",X"4E",X"12",X"57",X"12",X"59",X"12",X"63",X"12",
		X"6B",X"12",X"80",X"06",X"81",X"02",X"8F",X"13",X"92",X"0A",X"A0",X"03",X"A5",X"10",X"A8",X"07",
		X"B2",X"0F",X"B5",X"0F",X"C5",X"13",X"D4",X"09",X"E4",X"0F",X"E6",X"0C",X"F4",X"0C",X"04",X"10",
		X"06",X"0C",X"13",X"0C",X"20",X"06",X"21",X"03",X"22",X"10",X"23",X"19",X"28",X"10",X"2A",X"0A",
		X"3B",X"10",X"40",X"25",X"41",X"33",X"4A",X"1C",X"55",X"1C",X"65",X"1C",X"74",X"1C",X"82",X"0F",
		X"88",X"1C",X"95",X"0F",X"A5",X"1C",X"A8",X"30",X"B1",X"1C",X"B2",X"20",X"BE",X"0F",X"C0",X"06",
		X"C1",X"02",X"C2",X"1B",X"CA",X"10",X"E0",X"03",X"E6",X"0A",X"F0",X"17",X"03",X"08",X"12",X"18",
		X"13",X"09",X"40",X"1A",X"4A",X"0A",X"60",X"06",X"61",X"03",X"74",X"12",X"85",X"12",X"87",X"12",
		X"92",X"12",X"94",X"12",X"A9",X"12",X"AA",X"12",X"B4",X"10",X"BD",X"12",X"C3",X"12",X"CC",X"0F",
		X"D5",X"12",X"D7",X"12",X"E5",X"12",X"E7",X"12",X"F4",X"12",X"00",X"06",X"01",X"02",X"02",X"25",
		X"03",X"2C",X"0A",X"1C",X"17",X"1C",X"20",X"03",X"27",X"10",X"37",X"1C",X"48",X"1C",X"59",X"1C",
		X"6A",X"0A",X"79",X"1C",X"80",X"28",X"8D",X"0F",X"90",X"1C",X"91",X"20",X"A0",X"06",X"A1",X"03",
		X"AD",X"0C",X"B2",X"0F",X"BB",X"0C",X"CB",X"0C",X"D8",X"0F",X"E5",X"0F",X"E7",X"10",X"F1",X"0F",
		X"F9",X"0F",X"08",X"0C",X"0D",X"0F",X"16",X"0C",X"20",X"19",X"25",X"0F",X"28",X"09",X"36",X"10",
		X"40",X"06",X"41",X"02",X"42",X"25",X"4A",X"1C",X"5A",X"0F",X"60",X"03",X"61",X"2C",X"65",X"10",
		X"79",X"1C",X"88",X"1C",X"94",X"1C",X"A2",X"1C",X"AE",X"1C",X"BB",X"1C",X"BF",X"20",X"CA",X"0F",
		X"D0",X"28",X"DC",X"10",X"E0",X"06",X"E1",X"03",X"E8",X"0F",X"EA",X"10",X"EC",X"0A",X"F9",X"0F",
		X"08",X"13",X"0A",X"07",X"17",X"0F",X"1A",X"0A",X"2A",X"0C",X"37",X"10",X"3C",X"0C",X"43",X"02",
		X"80",X"06",X"00",X"06",X"20",X"03",X"28",X"10",X"34",X"0A",X"47",X"0C",X"55",X"0C",X"5A",X"0F",
		X"63",X"09",X"72",X"07",X"85",X"13",X"94",X"13",X"A0",X"06",X"A1",X"04",X"B3",X"14",X"BF",X"16",
		X"CD",X"16",X"DA",X"15",X"EC",X"16",X"EE",X"16",X"F8",X"16",X"F9",X"03",X"00",X"2B",X"20",X"23",
		X"40",X"86",X"4A",X"1C",X"50",X"28",X"65",X"1C",X"77",X"1C",X"7E",X"05",X"7F",X"20",X"80",X"33",
		X"C8",X"03",X"CF",X"30",X"E0",X"06",X"00",X"17",X"20",X"18",X"6A",X"0A",X"73",X"07",X"01",X"02",
		X"20",X"01",X"34",X"C0",X"3A",X"C2",X"48",X"20",X"54",X"C2",X"59",X"20",X"64",X"C2",X"69",X"E2",
		X"6D",X"C2",X"76",X"22",X"82",X"20",X"90",X"C0",X"96",X"C0",X"9C",X"C0",X"A2",X"C0",X"BE",X"C1",
		X"CB",X"C0",X"D8",X"20",X"E6",X"C2",X"F4",X"22",X"00",X"C2",X"05",X"FF",X"4D",X"00",X"4E",X"02",
		X"5E",X"22",X"77",X"22",X"8A",X"22",X"8B",X"FF",X"D8",X"00",X"E0",X"02",X"45",X"22",X"55",X"C2",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"46",X"E0",X"35",X"FB",X"78",X"32",X"13",X"E5",X"FE",X"05",X"CA",X"D2",X"27",X"A7",X"C2",
		X"5E",X"28",X"CD",X"FA",X"29",X"3E",X"1E",X"CD",X"75",X"0D",X"21",X"0F",X"E5",X"36",X"00",X"23",
		X"34",X"CD",X"48",X"29",X"CD",X"E8",X"05",X"21",X"24",X"2C",X"CD",X"00",X"03",X"CD",X"BA",X"28",
		X"21",X"0C",X"2C",X"CD",X"00",X"03",X"3A",X"13",X"E5",X"17",X"17",X"17",X"17",X"26",X"00",X"E6",
		X"F0",X"6F",X"20",X"01",X"24",X"22",X"98",X"E0",X"CD",X"71",X"29",X"2A",X"96",X"E0",X"56",X"2B",
		X"5E",X"2A",X"11",X"E5",X"A7",X"ED",X"52",X"30",X"0E",X"19",X"EB",X"2A",X"96",X"E0",X"72",X"2B",
		X"73",X"21",X"39",X"2C",X"CD",X"4E",X"03",X"2A",X"94",X"E0",X"ED",X"5B",X"11",X"E5",X"7D",X"D6",
		X"01",X"27",X"6F",X"30",X"01",X"25",X"22",X"94",X"E0",X"A7",X"ED",X"52",X"38",X"50",X"CD",X"68",
		X"29",X"2A",X"98",X"E0",X"7D",X"C6",X"01",X"27",X"6F",X"30",X"01",X"24",X"22",X"98",X"E0",X"CD",
		X"71",X"29",X"3E",X"10",X"CD",X"75",X"0D",X"3E",X"0C",X"CD",X"EA",X"05",X"18",X"C9",X"3E",X"1D",
		X"CD",X"75",X"0D",X"CD",X"D6",X"29",X"CD",X"12",X"0D",X"CD",X"48",X"29",X"3E",X"30",X"CD",X"EA",
		X"05",X"CD",X"BA",X"28",X"38",X"0D",X"21",X"E4",X"2B",X"CD",X"4E",X"03",X"3A",X"F9",X"E0",X"3C",
		X"C3",X"F9",X"27",X"21",X"F9",X"2B",X"CD",X"4E",X"03",X"CD",X"E8",X"05",X"18",X"0E",X"CD",X"E8",
		X"05",X"11",X"01",X"E5",X"21",X"98",X"E0",X"06",X"02",X"CD",X"36",X"06",X"21",X"00",X"00",X"22",
		X"11",X"E5",X"21",X"13",X"E5",X"7E",X"A7",X"C2",X"B7",X"0B",X"36",X"05",X"21",X"A2",X"23",X"22",
		X"16",X"E5",X"3E",X"1A",X"32",X"0E",X"E5",X"C3",X"B7",X"0B",X"CD",X"E8",X"05",X"CD",X"5A",X"29",
		X"3A",X"10",X"E5",X"D6",X"02",X"28",X"07",X"3E",X"0A",X"FA",X"CE",X"28",X"3E",X"05",X"5F",X"3A",
		X"13",X"E5",X"01",X"80",X"00",X"FE",X"08",X"30",X"09",X"01",X"00",X"01",X"FE",X"03",X"30",X"02",
		X"0E",X"20",X"ED",X"43",X"94",X"E0",X"83",X"87",X"5F",X"FE",X"0A",X"20",X"09",X"3A",X"10",X"E5",
		X"FE",X"03",X"28",X"02",X"1E",X"14",X"16",X"00",X"21",X"0C",X"E0",X"19",X"7E",X"23",X"22",X"96",
		X"E0",X"B6",X"20",X"03",X"70",X"2B",X"71",X"21",X"79",X"2B",X"CD",X"4E",X"03",X"CD",X"81",X"29",
		X"A7",X"20",X"02",X"3E",X"1A",X"C6",X"40",X"1B",X"1B",X"12",X"21",X"94",X"2B",X"CD",X"4E",X"03",
		X"21",X"12",X"E5",X"13",X"CD",X"9A",X"03",X"21",X"B0",X"2B",X"CD",X"4E",X"03",X"CD",X"68",X"29",
		X"21",X"CC",X"2B",X"CD",X"4E",X"03",X"2A",X"96",X"E0",X"13",X"CD",X"9A",X"03",X"2A",X"94",X"E0",
		X"ED",X"5B",X"11",X"E5",X"A7",X"ED",X"52",X"C9",X"21",X"00",X"E1",X"01",X"A4",X"00",X"CD",X"FA",
		X"05",X"01",X"20",X"02",X"21",X"E0",X"80",X"C3",X"FA",X"05",X"21",X"00",X"E1",X"01",X"C6",X"00",
		X"CD",X"FA",X"05",X"01",X"20",X"03",X"18",X"EC",X"11",X"D9",X"81",X"21",X"95",X"E0",X"C3",X"9A",
		X"03",X"21",X"99",X"E0",X"11",X"97",X"82",X"CD",X"93",X"03",X"EB",X"36",X"30",X"23",X"36",X"30",
		X"C9",X"3A",X"0E",X"E5",X"FE",X"1A",X"D8",X"D6",X"1A",X"C9",X"21",X"CC",X"80",X"11",X"CC",X"84",
		X"01",X"02",X"10",X"CD",X"E7",X"03",X"79",X"36",X"21",X"12",X"23",X"13",X"10",X"F9",X"21",X"CC",
		X"80",X"06",X"05",X"34",X"23",X"23",X"23",X"10",X"FA",X"36",X"1B",X"CD",X"81",X"29",X"21",X"CC",
		X"80",X"06",X"05",X"FE",X"05",X"38",X"0C",X"16",X"03",X"36",X"29",X"23",X"15",X"20",X"FA",X"D6",
		X"05",X"10",X"F0",X"57",X"87",X"87",X"82",X"5F",X"FE",X"08",X"38",X"10",X"28",X"01",X"3D",X"36",
		X"29",X"23",X"D6",X"08",X"18",X"F2",X"2A",X"F4",X"E0",X"3A",X"F6",X"E0",X"3C",X"57",X"C6",X"21",
		X"CB",X"66",X"28",X"07",X"D6",X"06",X"FE",X"20",X"20",X"01",X"3D",X"77",X"7A",X"FE",X"08",X"38",
		X"02",X"AF",X"2C",X"32",X"F6",X"E0",X"22",X"F4",X"E0",X"C9",X"21",X"CC",X"80",X"06",X"0F",X"36",
		X"29",X"23",X"10",X"FB",X"36",X"1F",X"3E",X"5A",X"32",X"52",X"80",X"C9",X"00",X"00",X"00",X"20",
		X"00",X"00",X"50",X"00",X"00",X"80",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",
		X"00",X"00",X"05",X"00",X"00",X"08",X"00",X"00",X"10",X"00",X"08",X"81",X"08",X"54",X"4F",X"20",
		X"43",X"4F",X"55",X"4E",X"54",X"49",X"4E",X"55",X"45",X"20",X"47",X"41",X"4D",X"45",X"22",X"2D",
		X"82",X"08",X"54",X"49",X"4D",X"45",X"21",X"46",X"81",X"08",X"42",X"45",X"47",X"49",X"4E",X"4E",
		X"45",X"52",X"20",X"43",X"4F",X"55",X"52",X"53",X"45",X"20",X"47",X"4F",X"20",X"5B",X"21",X"46",
		X"81",X"00",X"43",X"48",X"41",X"4D",X"50",X"49",X"4F",X"4E",X"20",X"43",X"4F",X"55",X"52",X"53",
		X"45",X"20",X"31",X"20",X"47",X"4F",X"20",X"5B",X"21",X"4C",X"82",X"00",X"46",X"52",X"45",X"45",
		X"20",X"50",X"4C",X"41",X"59",X"21",X"EA",X"81",X"00",X"4F",X"4E",X"4C",X"59",X"20",X"31",X"20",
		X"50",X"4C",X"41",X"59",X"45",X"52",X"21",X"EA",X"81",X"00",X"31",X"20",X"4F",X"52",X"20",X"32",
		X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"53",X"21",X"06",X"82",X"00",X"50",X"49",X"43",X"54",
		X"55",X"52",X"45",X"20",X"4E",X"55",X"4D",X"42",X"45",X"52",X"20",X"53",X"45",X"54",X"22",X"4A",
		X"82",X"00",X"4E",X"45",X"58",X"54",X"20",X"31",X"50",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"21",X"6A",X"81",X"00",X"20",X"50",X"55",X"53",X"48",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"20",X"21",X"D4",X"83",X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"21",X"88",X"81",X"00",
		X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"20",X"21",X"0C",X"82",X"00",X"47",X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"21",X"2B",
		X"80",X"02",X"04",X"25",X"0F",X"14",X"05",X"22",X"41",X"80",X"01",X"0C",X"0D",X"25",X"06",X"00",
		X"22",X"49",X"80",X"09",X"3F",X"22",X"4B",X"80",X"02",X"06",X"50",X"4F",X"49",X"4E",X"54",X"25",
		X"04",X"00",X"12",X"25",X"05",X"00",X"07",X"22",X"6B",X"80",X"02",X"06",X"25",X"09",X"00",X"12",
		X"25",X"05",X"00",X"07",X"22",X"8B",X"80",X"02",X"06",X"0E",X"0F",X"10",X"11",X"25",X"05",X"00",
		X"12",X"25",X"05",X"00",X"07",X"22",X"AB",X"80",X"02",X"08",X"16",X"15",X"15",X"17",X"15",X"15",
		X"18",X"15",X"15",X"19",X"15",X"15",X"1A",X"15",X"15",X"09",X"22",X"81",X"80",X"01",X"31",X"50",
		X"3F",X"21",X"A1",X"80",X"01",X"32",X"50",X"3F",X"21",X"25",X"81",X"01",X"54",X"49",X"4D",X"45",
		X"20",X"54",X"4F",X"20",X"52",X"45",X"41",X"43",X"48",X"20",X"50",X"4F",X"49",X"4E",X"54",X"20",
		X"5E",X"00",X"5E",X"21",X"84",X"81",X"00",X"59",X"4F",X"55",X"52",X"20",X"54",X"49",X"4D",X"45",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"22",X"97",X"81",X"01",X"5D",X"21",
		X"C4",X"81",X"00",X"54",X"48",X"45",X"20",X"41",X"56",X"45",X"52",X"41",X"47",X"45",X"20",X"54",
		X"49",X"4D",X"45",X"20",X"20",X"20",X"22",X"D7",X"81",X"01",X"5D",X"21",X"04",X"82",X"01",X"54",
		X"4F",X"50",X"20",X"52",X"45",X"43",X"4F",X"52",X"44",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"5D",X"21",X"85",X"82",X"00",X"47",X"4F",X"4F",X"44",X"20",X"42",X"4F",X"4E",X"55",
		X"53",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"21",X"67",X"82",X"00",X"53",X"4F",X"52",X"52",
		X"59",X"20",X"4E",X"4F",X"20",X"42",X"4F",X"4E",X"55",X"53",X"5B",X"21",X"65",X"82",X"01",X"53",
		X"50",X"45",X"43",X"49",X"41",X"4C",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"21",X"25",X"81",X"00",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",X"55",X"4C",
		X"41",X"54",X"49",X"4F",X"4E",X"53",X"20",X"5B",X"21",X"E5",X"82",X"01",X"59",X"4F",X"55",X"20",
		X"48",X"41",X"56",X"45",X"20",X"42",X"52",X"4F",X"4B",X"45",X"4E",X"20",X"41",X"20",X"52",X"45",
		X"43",X"4F",X"52",X"44",X"20",X"5B",X"21",X"6A",X"81",X"00",X"49",X"4E",X"53",X"45",X"52",X"54",
		X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"C7",X"81",X"00",X"31",X"20",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"20",X"20",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"C5",X"81",X"00",
		X"41",X"20",X"5F",X"20",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"20",X"20",X"31",
		X"20",X"43",X"4F",X"49",X"4E",X"20",X"21",X"C8",X"82",X"00",X"5C",X"31",X"39",X"38",X"32",X"20",
		X"49",X"52",X"45",X"4D",X"20",X"43",X"4F",X"52",X"50",X"2F",X"21",X"76",X"80",X"02",X"3A",X"3B",
		X"3C",X"3D",X"3E",X"21",X"F0",X"F0",X"ED",X"F0",X"F0",X"FB",X"FB",X"FB",X"F0",X"E8",X"F0",X"F0",
		X"F0",X"EE",X"F0",X"F0",X"F0",X"F0",X"E0",X"F0",X"F0",X"FB",X"FB",X"FB",X"F0",X"F0",X"F0",X"F2",
		X"F2",X"F0",X"F0",X"F0",X"E9",X"F2",X"EF",X"E3",X"D2",X"FC",X"FD",X"FE",X"E0",X"D4",X"D3",X"EB",
		X"FF",X"D5",X"F1",X"E5",X"E2",X"D0",X"D6",X"E6",X"D7",X"F0",X"E1",X"D8",X"F9",X"FB",X"F0",X"F2",
		X"D9",X"EC",X"FC",X"D1",X"34",X"32",X"32",X"43",X"34",X"23",X"32",X"11",X"23",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"12",X"12",X"12",X"24",X"77",X"21",X"10",X"56",X"21",X"10",X"34",X"21",
		X"23",X"23",X"21",X"31",X"22",X"21",X"11",X"00",X"77",X"77",X"66",X"65",X"55",X"44",X"43",X"33",
		X"43",X"33",X"21",X"31",X"00",X"9A",X"51",X"98",X"8D",X"5F",X"B6",X"30",X"D2",X"06",X"E3",X"E3",
		X"EF",X"C7",X"F7",X"B0",X"FC",X"9E",X"00",X"8E",X"03",X"82",X"06",X"77",X"07",X"6E",X"08",X"66",
		X"09",X"5F",X"0A",X"59",X"03",X"48",X"81",X"B0",X"B1",X"B2",X"B3",X"B4",X"02",X"B5",X"B6",X"B7",
		X"B8",X"02",X"B9",X"BA",X"BB",X"BC",X"BD",X"02",X"BE",X"BF",X"C0",X"C1",X"C2",X"02",X"C3",X"C4",
		X"C5",X"C6",X"BD",X"02",X"03",X"6D",X"81",X"C7",X"C8",X"C9",X"CA",X"02",X"CB",X"BF",X"CC",X"02",
		X"CD",X"BC",X"CE",X"CF",X"02",X"D0",X"D1",X"D2",X"CA",X"02",X"D3",X"D4",X"D5",X"C2",X"02",X"D6",
		X"D7",X"BC",X"BD",X"02",X"D8",X"C0",X"C1",X"C2",X"02",X"D9",X"BC",X"C5",X"DA",X"02",X"DB",X"C1",
		X"DC",X"02",X"03",X"06",X"82",X"B0",X"B1",X"B2",X"B3",X"B4",X"02",X"DD",X"DE",X"DF",X"B8",X"02",
		X"E0",X"E1",X"E2",X"02",X"E3",X"E4",X"E5",X"02",X"00",X"E6",X"B2",X"E7",X"E8",X"02",X"00",X"E9",
		X"EA",X"EB",X"EC",X"02",X"00",X"ED",X"EE",X"EF",X"B4",X"02",X"00",X"F0",X"F1",X"F2",X"02",X"F3",
		X"F4",X"F5",X"BF",X"02",X"F7",X"F8",X"F9",X"B0",X"FA",X"02",X"00",X"B2",X"B3",X"FB",X"FC",X"02",
		X"00",X"FD",X"B8",X"02",X"00",X"FE",X"BC",X"CE",X"CF",X"02",X"00",X"D0",X"D1",X"D2",X"CA",X"02",
		X"00",X"D3",X"D4",X"D5",X"C2",X"02",X"00",X"D6",X"D7",X"BC",X"BD",X"02",X"C5",X"BF",X"C0",X"FF",
		X"EC",X"02",X"C3",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"19",X"2F",X"08",X"02",X"18",X"2F",X"08",X"02",X"15",X"38",X"0D",X"04",X"15",X"38",X"0D",X"04",
		X"15",X"42",X"10",X"04",X"15",X"33",X"10",X"00",X"01",X"00",X"0E",X"04",X"09",X"00",X"24",X"04",
		X"0D",X"00",X"24",X"04",X"11",X"01",X"08",X"06",X"17",X"01",X"08",X"06",X"1D",X"01",X"08",X"06",
		X"23",X"01",X"0A",X"02",X"25",X"01",X"0A",X"02",X"27",X"01",X"0C",X"01",X"28",X"01",X"1C",X"01",
		X"29",X"01",X"1C",X"01",X"2A",X"01",X"1C",X"01",X"2B",X"01",X"1C",X"01",X"2C",X"01",X"1C",X"01",
		X"2D",X"04",X"00",X"01",X"2E",X"04",X"00",X"01",X"2F",X"04",X"00",X"01",X"30",X"04",X"00",X"01",
		X"31",X"04",X"00",X"01",X"31",X"84",X"00",X"01",X"31",X"C4",X"00",X"01",X"31",X"44",X"00",X"01",
		X"32",X"04",X"00",X"01",X"33",X"04",X"00",X"01",X"34",X"04",X"00",X"01",X"33",X"C4",X"00",X"01",
		X"34",X"C4",X"00",X"01",X"36",X"04",X"00",X"01",X"36",X"84",X"00",X"01",X"37",X"04",X"00",X"01",
		X"36",X"C4",X"00",X"01",X"36",X"44",X"00",X"01",X"37",X"C4",X"00",X"01",X"38",X"09",X"00",X"01",
		X"39",X"00",X"00",X"01",X"3A",X"09",X"02",X"02",X"05",X"00",X"2C",X"01",X"3D",X"0A",X"28",X"01",
		X"3E",X"01",X"00",X"01",X"3F",X"01",X"00",X"01",X"40",X"01",X"00",X"01",X"41",X"01",X"00",X"01",
		X"42",X"07",X"1A",X"80",X"45",X"07",X"1A",X"80",X"46",X"07",X"1A",X"80",X"47",X"07",X"1A",X"80",
		X"47",X"47",X"1A",X"80",X"46",X"47",X"1A",X"80",X"45",X"47",X"1A",X"80",X"43",X"07",X"1A",X"01",
		X"44",X"07",X"1A",X"01",X"43",X"87",X"1A",X"01",X"44",X"47",X"1A",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"48",X"01",X"1A",X"80",X"49",X"01",X"1A",X"80",X"4A",X"01",X"1A",X"80",
		X"35",X"0A",X"2A",X"80",X"4B",X"01",X"1A",X"80",X"4C",X"01",X"1A",X"80",X"4D",X"01",X"1A",X"80",
		X"4E",X"01",X"00",X"C0",X"4F",X"01",X"10",X"C0",X"53",X"01",X"10",X"C0",X"57",X"01",X"10",X"C0",
		X"5B",X"01",X"12",X"C0",X"61",X"03",X"1E",X"C0",X"62",X"03",X"1E",X"C0",X"63",X"03",X"1E",X"C0",
		X"64",X"03",X"14",X"C0",X"68",X"03",X"14",X"C0",X"6C",X"03",X"16",X"C0",X"6E",X"03",X"16",X"C0",
		X"78",X"08",X"22",X"02",X"70",X"02",X"04",X"04",X"73",X"02",X"06",X"04",X"74",X"02",X"18",X"04",
		X"75",X"02",X"20",X"04",X"7A",X"01",X"1A",X"80",X"4B",X"41",X"1A",X"80",X"4C",X"41",X"1A",X"80",
		X"7B",X"09",X"26",X"02",X"07",X"00",X"2C",X"01",X"7D",X"0E",X"2E",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A3",
		X"01",X"02",X"02",X"03",X"03",X"04",X"04",X"05",X"60",X"01",X"58",X"01",X"50",X"01",X"48",X"01",
		X"40",X"01",X"38",X"01",X"39",X"10",X"39",X"20",X"39",X"30",X"39",X"48",X"39",X"60",X"39",X"70",
		X"39",X"80",X"39",X"98",X"39",X"B0",X"39",X"D0",X"B4",X"38",X"FF",X"58",X"8E",X"28",X"B4",X"38",
		X"00",X"19",X"24",X"2C",X"33",X"39",X"3E",X"43",X"48",X"4C",X"50",X"54",X"58",X"5B",X"5F",X"62",
		X"65",X"68",X"6B",X"6E",X"71",X"74",X"77",X"79",X"7C",X"7E",X"50",X"5E",X"6B",X"87",X"87",X"A2",
		X"A2",X"A3",X"02",X"00",X"A4",X"A5",X"02",X"00",X"A6",X"A7",X"02",X"A8",X"A9",X"01",X"AA",X"02",
		X"AB",X"AC",X"AD",X"02",X"00",X"AE",X"AF",X"02",X"B0",X"B1",X"01",X"B2",X"B3",X"B4",X"02",X"00",
		X"B5",X"B6",X"B7",X"02",X"00",X"00",X"00",X"B8",X"B9",X"02",X"00",X"00",X"00",X"BA",X"02",X"00",
		X"BB",X"BC",X"BD",X"02",X"BE",X"BF",X"01",X"C0",X"C1",X"02",X"00",X"C2",X"C3",X"C4",X"02",X"00",
		X"00",X"00",X"C5",X"C6",X"02",X"00",X"00",X"00",X"C7",X"C8",X"02",X"00",X"C9",X"CA",X"CB",X"02",
		X"CC",X"01",X"DA",X"DB",X"DC",X"02",X"00",X"00",X"F0",X"03",X"00",X"00",X"F0",X"02",X"00",X"00",
		X"F0",X"02",X"DD",X"DE",X"DF",X"01",X"0F",X"04",X"05",X"0F",X"24",X"27",X"0F",X"43",X"48",X"11",
		X"48",X"4E",X"12",X"4E",X"53",X"10",X"63",X"68",X"13",X"68",X"6C",X"0F",X"6C",X"6D",X"14",X"6D",
		X"6E",X"12",X"6E",X"74",X"10",X"89",X"8E",X"FF",X"0C",X"03",X"03",X"03",X"02",X"01",X"FF",X"3B",
		X"FF",X"70",X"FC",X"24",X"B9",X"FF",X"10",X"FC",X"24",X"3B",X"01",X"A0",X"FC",X"53",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0A",X"0D",X"0F",X"11",X"13",X"15",X"16",X"18",X"19",X"1A",X"1B",X"1D",X"1E",X"1F",X"20",
		X"21",X"22",X"23",X"24",X"25",X"26",X"27",X"28",X"28",X"28",X"28",X"28",X"FF",X"1F",X"01",X"1C",
		X"04",X"0C",X"00",X"24",X"02",X"1D",X"05",X"20",X"08",X"0C",X"04",X"34",X"05",X"21",X"06",X"07",
		X"07",X"0C",X"0C",X"14",X"05",X"1E",X"08",X"1E",X"0F",X"0C",X"12",X"34",X"02",X"1B",X"03",X"1A",
		X"06",X"10",X"21",X"42",X"02",X"1D",X"04",X"1D",X"08",X"0F",X"27",X"42",X"05",X"20",X"06",X"20",
		X"0B",X"0C",X"2F",X"42",X"09",X"16",X"02",X"22",X"06",X"1C",X"3A",X"4E",X"0E",X"19",X"03",X"26",
		X"07",X"1C",X"40",X"4E",X"12",X"1D",X"05",X"2A",X"0A",X"1C",X"47",X"4E",X"05",X"20",X"05",X"26",
		X"08",X"0C",X"51",X"45",X"05",X"19",X"05",X"1F",X"11",X"0C",X"58",X"7F",X"08",X"1E",X"04",X"1E",
		X"09",X"0C",X"69",X"00",X"00",X"1B",X"16",X"1C",X"17",X"1A",X"72",X"20",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"04",X"03",X"01",X"01",X"03",X"04",X"06",X"07",X"08",X"07",X"05",X"02",X"04",X"06",X"08",
		X"09",X"0B",X"01",X"03",X"04",X"06",X"07",X"09",X"0A",X"0C",X"0D",X"0C",X"0A",X"08",X"07",X"05",
		X"03",X"01",X"02",X"04",X"05",X"04",X"02",X"01",X"03",X"05",X"06",X"08",X"07",X"05",X"03",X"02",
		X"04",X"06",X"08",X"0A",X"0B",X"0D",X"0B",X"09",X"07",X"05",X"01",X"02",X"03",X"02",X"02",X"01",
		X"04",X"06",X"07",X"08",X"06",X"04",X"01",X"02",X"04",X"06",X"08",X"0A",X"0C",X"0B",X"0A",X"05",
		X"02",X"03",X"07",X"09",X"0A",X"0C",X"0B",X"09",X"03",X"03",X"07",X"09",X"09",X"0B",X"0A",X"0A",
		X"0A",X"09",X"08",X"08",X"07",X"06",X"06",X"04",X"04",X"02",X"04",X"05",X"07",X"08",X"07",X"05",
		X"03",X"00",X"02",X"02",X"02",X"02",X"02",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"F8",X"02",X"02",
		X"02",X"02",X"02",X"F8",X"F8",X"F8",X"F8",X"F8",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3E",X"FF",X"D3",X"C0",X"32",X"C5",X"E1",X"21",X"00",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",
		X"CF",X"00",X"ED",X"B0",X"3E",X"01",X"57",X"01",X"00",X"08",X"21",X"00",X"E0",X"7A",X"77",X"5E",
		X"BB",X"C2",X"BB",X"34",X"23",X"0B",X"79",X"B0",X"20",X"F3",X"7A",X"07",X"30",X"E8",X"16",X"55",
		X"7A",X"01",X"00",X"08",X"21",X"00",X"E0",X"77",X"23",X"3C",X"5F",X"0B",X"79",X"B0",X"28",X"09",
		X"7B",X"FE",X"AB",X"20",X"F2",X"3E",X"55",X"18",X"EE",X"7A",X"01",X"00",X"08",X"21",X"00",X"E0",
		X"BE",X"20",X"19",X"23",X"3C",X"5F",X"0B",X"79",X"B0",X"28",X"09",X"7B",X"FE",X"AB",X"20",X"F0",
		X"3E",X"55",X"18",X"EC",X"14",X"7A",X"FE",X"AB",X"20",X"C6",X"18",X"09",X"5E",X"57",X"AF",X"C3",
		X"BB",X"34",X"7A",X"18",X"DE",X"31",X"00",X"E8",X"3E",X"01",X"57",X"01",X"00",X"08",X"21",X"00",
		X"80",X"7A",X"77",X"5E",X"BB",X"28",X"08",X"CD",X"3B",X"35",X"CB",X"4F",X"CA",X"F5",X"33",X"23",
		X"0B",X"79",X"B0",X"20",X"EC",X"7A",X"07",X"30",X"E1",X"16",X"55",X"7A",X"01",X"00",X"08",X"21",
		X"00",X"80",X"77",X"23",X"3C",X"5F",X"0B",X"79",X"B0",X"28",X"09",X"7B",X"FE",X"AB",X"20",X"F2",
		X"3E",X"55",X"18",X"EE",X"7A",X"01",X"00",X"08",X"21",X"00",X"80",X"BE",X"20",X"19",X"23",X"3C",
		X"5F",X"0B",X"79",X"B0",X"28",X"09",X"7B",X"FE",X"AB",X"20",X"F0",X"3E",X"55",X"18",X"EC",X"14",
		X"7A",X"FE",X"AB",X"20",X"C6",X"18",X"0D",X"5E",X"57",X"CD",X"37",X"35",X"CB",X"4F",X"CA",X"F5",
		X"33",X"7A",X"18",X"DA",X"DD",X"21",X"EB",X"33",X"C3",X"B1",X"35",X"21",X"66",X"3A",X"DD",X"21",
		X"F5",X"33",X"C3",X"65",X"34",X"21",X"00",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",X"CF",X"00",
		X"ED",X"B0",X"21",X"00",X"00",X"AF",X"32",X"00",X"E7",X"06",X"00",X"0E",X"10",X"AF",X"AE",X"23",
		X"10",X"FC",X"0D",X"20",X"F9",X"E5",X"CD",X"35",X"34",X"E1",X"3A",X"00",X"E7",X"3C",X"FE",X"04",
		X"20",X"E4",X"AF",X"D3",X"1C",X"FB",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"F9",X"3E",X"03",X"32",
		X"01",X"E7",X"C3",X"CD",X"35",X"F5",X"FE",X"FF",X"28",X"02",X"0E",X"08",X"21",X"86",X"3A",X"09",
		X"EB",X"3A",X"00",X"E7",X"0F",X"0F",X"4F",X"21",X"C4",X"80",X"09",X"E5",X"EB",X"0E",X"08",X"ED",
		X"B0",X"13",X"13",X"D5",X"FD",X"E1",X"DD",X"E1",X"F1",X"CD",X"9A",X"34",X"3A",X"00",X"E7",X"C6",
		X"30",X"DD",X"77",X"03",X"C9",X"7E",X"23",X"FE",X"00",X"28",X"0B",X"5E",X"23",X"56",X"23",X"4F",
		X"06",X"00",X"ED",X"B0",X"18",X"EF",X"DD",X"E9",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C6",X"30",
		X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"00",X"DD",X"E9",X"E6",X"0F",X"C6",X"30",X"FE",
		X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"01",X"DD",X"E9",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"00",X"F1",X"E6",X"0F",X"C6",
		X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"FD",X"77",X"01",X"C9",X"08",X"D9",X"DD",X"21",X"C4",
		X"34",X"C3",X"B1",X"35",X"21",X"72",X"3A",X"DD",X"21",X"CE",X"34",X"C3",X"65",X"34",X"D9",X"FD",
		X"21",X"8F",X"80",X"DD",X"21",X"DB",X"34",X"7C",X"C3",X"78",X"34",X"DD",X"21",X"E3",X"34",X"7C",
		X"C3",X"8B",X"34",X"FD",X"23",X"FD",X"23",X"DD",X"21",X"EF",X"34",X"7D",X"C3",X"78",X"34",X"DD",
		X"21",X"F7",X"34",X"7D",X"C3",X"8B",X"34",X"FD",X"21",X"95",X"80",X"DD",X"21",X"03",X"35",X"7A",
		X"C3",X"78",X"34",X"DD",X"21",X"0B",X"35",X"7A",X"C3",X"8B",X"34",X"FD",X"21",X"99",X"80",X"DD",
		X"21",X"17",X"35",X"7B",X"C3",X"78",X"34",X"7B",X"DD",X"21",X"1F",X"35",X"C3",X"8B",X"34",X"3A",
		X"00",X"D0",X"CB",X"47",X"CA",X"2F",X"35",X"CB",X"4F",X"20",X"F4",X"08",X"C3",X"F5",X"33",X"08",
		X"B7",X"CA",X"72",X"33",X"C3",X"24",X"33",X"E5",X"D9",X"18",X"09",X"E5",X"D9",X"DD",X"21",X"44",
		X"35",X"C3",X"B1",X"35",X"21",X"00",X"80",X"11",X"00",X"E0",X"01",X"A0",X"04",X"ED",X"B0",X"21",
		X"00",X"80",X"36",X"00",X"54",X"5D",X"13",X"01",X"9F",X"04",X"ED",X"B0",X"21",X"72",X"3A",X"DD",
		X"21",X"66",X"35",X"C3",X"65",X"34",X"D9",X"FD",X"21",X"8F",X"80",X"7C",X"CD",X"9A",X"34",X"FD",
		X"23",X"FD",X"23",X"7D",X"CD",X"9A",X"34",X"FD",X"21",X"95",X"80",X"7A",X"CD",X"9A",X"34",X"FD",
		X"21",X"99",X"80",X"7B",X"CD",X"9A",X"34",X"E1",X"3A",X"00",X"D0",X"CB",X"47",X"28",X"06",X"CB",
		X"4F",X"28",X"10",X"18",X"F3",X"D9",X"21",X"00",X"E0",X"11",X"00",X"80",X"01",X"A0",X"04",X"ED",
		X"B0",X"D9",X"C9",X"21",X"A0",X"84",X"36",X"00",X"54",X"5D",X"13",X"01",X"5F",X"03",X"ED",X"B0",
		X"C9",X"21",X"00",X"84",X"01",X"FF",X"03",X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"21",X"00",
		X"80",X"01",X"FF",X"03",X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"DD",X"E9",X"CD",X"AD",X"38",
		X"21",X"BF",X"3E",X"CD",X"08",X"39",X"3A",X"01",X"E7",X"06",X"02",X"CD",X"1C",X"39",X"3A",X"00",
		X"D0",X"CB",X"47",X"20",X"14",X"3A",X"01",X"E7",X"07",X"4F",X"06",X"00",X"DD",X"21",X"96",X"3A",
		X"DD",X"09",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E9",X"DD",X"21",X"02",X"E7",X"CD",X"DD",X"38",
		X"47",X"E6",X"55",X"FE",X"55",X"28",X"09",X"78",X"E6",X"AA",X"FE",X"AA",X"28",X"13",X"18",X"CE",
		X"DD",X"36",X"00",X"55",X"DD",X"36",X"01",X"08",X"DD",X"36",X"02",X"01",X"CD",X"32",X"36",X"18",
		X"BD",X"DD",X"36",X"00",X"AA",X"DD",X"36",X"01",X"03",X"DD",X"36",X"02",X"FF",X"CD",X"32",X"36",
		X"18",X"AC",X"DD",X"56",X"00",X"1E",X"02",X"CD",X"C8",X"38",X"28",X"0E",X"CD",X"4E",X"36",X"DD",
		X"56",X"00",X"1E",X"01",X"CD",X"C8",X"38",X"20",X"F3",X"C9",X"CD",X"4E",X"36",X"C9",X"3A",X"01",
		X"E7",X"DD",X"BE",X"01",X"C8",X"06",X"00",X"CD",X"1C",X"39",X"DD",X"86",X"02",X"32",X"01",X"E7",
		X"06",X"02",X"CD",X"1C",X"39",X"C9",X"CD",X"AD",X"38",X"21",X"10",X"3B",X"CD",X"08",X"39",X"3A",
		X"03",X"D0",X"21",X"CB",X"80",X"CD",X"B2",X"36",X"3A",X"04",X"D0",X"21",X"0B",X"81",X"CD",X"B2",
		X"36",X"DD",X"21",X"AC",X"3A",X"FD",X"21",X"A8",X"3A",X"3A",X"03",X"D0",X"EE",X"FF",X"06",X"02",
		X"CD",X"C6",X"36",X"DD",X"21",X"F8",X"3A",X"FD",X"21",X"F4",X"3A",X"3A",X"04",X"D0",X"EE",X"FF",
		X"06",X"01",X"CD",X"C5",X"36",X"CD",X"EC",X"36",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"C0",X"C3",
		X"CD",X"35",X"EE",X"FF",X"06",X"08",X"0F",X"38",X"04",X"36",X"30",X"18",X"02",X"36",X"31",X"23",
		X"23",X"10",X"F3",X"C9",X"0F",X"0F",X"4F",X"C5",X"DD",X"A6",X"00",X"DD",X"86",X"01",X"DD",X"23",
		X"DD",X"23",X"4F",X"06",X"00",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"09",X"4E",X"FD",X"6E",X"02",
		X"FD",X"66",X"03",X"09",X"CD",X"11",X"39",X"C1",X"79",X"10",X"D9",X"C9",X"3A",X"04",X"D0",X"CB",
		X"57",X"CA",X"06",X"37",X"21",X"77",X"3B",X"CD",X"08",X"39",X"DD",X"21",X"99",X"3B",X"FD",X"21",
		X"9B",X"3B",X"06",X"01",X"18",X"10",X"21",X"7F",X"3C",X"CD",X"08",X"39",X"DD",X"21",X"92",X"3C",
		X"FD",X"21",X"96",X"3C",X"06",X"02",X"3A",X"03",X"D0",X"EE",X"FF",X"0F",X"0F",X"CD",X"C4",X"36",
		X"C9",X"AF",X"32",X"0F",X"E7",X"67",X"6F",X"22",X"0D",X"E7",X"CD",X"AD",X"38",X"21",X"22",X"3D",
		X"CD",X"08",X"39",X"3A",X"00",X"D0",X"21",X"CB",X"80",X"CD",X"B2",X"36",X"3A",X"01",X"D0",X"21",
		X"0B",X"81",X"CD",X"B2",X"36",X"3A",X"02",X"D0",X"21",X"4B",X"81",X"CD",X"B2",X"36",X"CD",X"8C",
		X"37",X"3A",X"0D",X"E7",X"21",X"8C",X"81",X"CD",X"7A",X"37",X"23",X"3A",X"0E",X"E7",X"CD",X"7A",
		X"37",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"CB",X"3A",X"01",X"D0",X"CB",X"4F",X"20",X"C4",X"CD",
		X"AD",X"38",X"3E",X"01",X"CD",X"3C",X"39",X"C3",X"CD",X"35",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",
		X"0F",X"C6",X"30",X"77",X"23",X"F1",X"E6",X"0F",X"C6",X"30",X"77",X"C9",X"21",X"0F",X"E7",X"3A",
		X"4E",X"E0",X"E6",X"C0",X"BE",X"C8",X"32",X"0F",X"E7",X"3A",X"0E",X"E7",X"C6",X"01",X"27",X"32",
		X"0E",X"E7",X"D0",X"3A",X"0D",X"E7",X"C6",X"01",X"27",X"32",X"0D",X"E7",X"C9",X"2A",X"53",X"3D",
		X"22",X"06",X"E7",X"21",X"68",X"3D",X"FD",X"21",X"57",X"3D",X"CD",X"C0",X"37",X"C3",X"CD",X"35",
		X"FD",X"22",X"0B",X"E7",X"E5",X"CD",X"AD",X"38",X"E1",X"CD",X"08",X"39",X"DD",X"21",X"08",X"E7",
		X"3E",X"01",X"32",X"05",X"E7",X"06",X"02",X"CD",X"23",X"39",X"3E",X"01",X"0E",X"40",X"CD",X"3E",
		X"39",X"CD",X"72",X"38",X"CD",X"7D",X"38",X"3E",X"FF",X"32",X"11",X"E7",X"3A",X"00",X"D0",X"CB",
		X"4F",X"28",X"4A",X"CD",X"F2",X"38",X"E6",X"AA",X"FE",X"2A",X"28",X"13",X"CD",X"DD",X"38",X"47",
		X"E6",X"55",X"FE",X"55",X"28",X"11",X"78",X"E6",X"AA",X"FE",X"AA",X"28",X"1D",X"18",X"DD",X"CD",
		X"72",X"38",X"CD",X"7D",X"38",X"18",X"D5",X"DD",X"36",X"00",X"55",X"3A",X"06",X"E7",X"DD",X"77",
		X"01",X"DD",X"36",X"02",X"01",X"CD",X"4F",X"38",X"18",X"C2",X"DD",X"36",X"00",X"AA",X"3A",X"07",
		X"E7",X"DD",X"77",X"01",X"DD",X"36",X"02",X"FF",X"CD",X"4F",X"38",X"18",X"AF",X"CD",X"72",X"38",
		X"3E",X"01",X"0E",X"20",X"CD",X"3E",X"39",X"3A",X"00",X"D0",X"CB",X"4F",X"20",X"9E",X"C9",X"CD",
		X"72",X"38",X"DD",X"56",X"00",X"1E",X"02",X"CD",X"C8",X"38",X"28",X"0F",X"CD",X"95",X"38",X"DD",
		X"56",X"00",X"1E",X"01",X"CD",X"C8",X"38",X"20",X"F3",X"18",X"03",X"CD",X"95",X"38",X"CD",X"7D",
		X"38",X"C9",X"3E",X"00",X"32",X"00",X"D0",X"CB",X"FF",X"32",X"00",X"D0",X"C9",X"3A",X"05",X"E7",
		X"4F",X"06",X"00",X"FD",X"2A",X"0B",X"E7",X"FD",X"09",X"FD",X"7E",X"00",X"32",X"00",X"D0",X"CB",
		X"FF",X"32",X"00",X"D0",X"C9",X"3A",X"05",X"E7",X"DD",X"BE",X"01",X"C8",X"06",X"00",X"CD",X"23",
		X"39",X"DD",X"86",X"02",X"32",X"05",X"E7",X"06",X"02",X"CD",X"23",X"39",X"C9",X"21",X"00",X"80",
		X"01",X"FF",X"03",X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"21",X"00",X"84",X"01",X"FF",X"03",
		X"36",X"00",X"54",X"5D",X"13",X"ED",X"B0",X"C9",X"0E",X"00",X"06",X"0C",X"CD",X"E2",X"38",X"A2",
		X"C8",X"10",X"F9",X"0D",X"20",X"F4",X"1D",X"20",X"EF",X"3E",X"FF",X"A2",X"C9",X"CD",X"E2",X"38",
		X"18",X"1F",X"21",X"10",X"E7",X"3A",X"01",X"D0",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"EE",
		X"FF",X"C9",X"21",X"11",X"E7",X"3A",X"00",X"D0",X"1F",X"CB",X"16",X"1F",X"CB",X"16",X"7E",X"EE",
		X"FF",X"F5",X"AF",X"3D",X"20",X"FD",X"F1",X"C9",X"7E",X"FE",X"00",X"C8",X"CD",X"11",X"39",X"18",
		X"F7",X"4E",X"06",X"00",X"23",X"5E",X"23",X"56",X"23",X"ED",X"B0",X"C9",X"4F",X"D6",X"03",X"07",
		X"3C",X"18",X"01",X"4F",X"C5",X"0E",X"64",X"06",X"00",X"60",X"07",X"07",X"07",X"6F",X"29",X"29",
		X"09",X"EB",X"21",X"00",X"84",X"19",X"C1",X"70",X"23",X"70",X"79",X"C9",X"0E",X"00",X"06",X"00",
		X"10",X"FE",X"0D",X"20",X"F9",X"3D",X"20",X"F4",X"C9",X"C5",X"0E",X"00",X"06",X"00",X"10",X"FE",
		X"F5",X"3A",X"00",X"D0",X"CB",X"4F",X"28",X"09",X"F1",X"0D",X"20",X"F0",X"3D",X"20",X"EB",X"C1",
		X"C9",X"F1",X"C1",X"06",X"01",X"C9",X"CD",X"AD",X"38",X"11",X"00",X"E1",X"21",X"6D",X"3E",X"01",
		X"10",X"00",X"ED",X"B0",X"11",X"60",X"E1",X"21",X"7D",X"3E",X"01",X"10",X"00",X"ED",X"B0",X"3A",
		X"00",X"D0",X"CB",X"4F",X"20",X"F9",X"21",X"00",X"E1",X"36",X"00",X"54",X"5D",X"13",X"01",X"BF",
		X"00",X"ED",X"B0",X"C3",X"CD",X"35",X"3E",X"01",X"32",X"12",X"E7",X"AF",X"32",X"11",X"E7",X"18",
		X"2A",X"3A",X"00",X"D0",X"CB",X"4F",X"CA",X"CD",X"35",X"CD",X"F2",X"38",X"E6",X"AA",X"FE",X"2A",
		X"20",X"EF",X"3A",X"12",X"E7",X"3C",X"32",X"12",X"E7",X"FE",X"01",X"28",X"0E",X"FE",X"02",X"CA",
		X"E8",X"39",X"FE",X"03",X"CA",X"13",X"3A",X"D6",X"03",X"18",X"EB",X"CD",X"AD",X"38",X"21",X"1C",
		X"81",X"06",X"1A",X"3E",X"5A",X"77",X"2B",X"3D",X"10",X"FB",X"21",X"0C",X"82",X"06",X"0A",X"3E",
		X"39",X"77",X"2B",X"3D",X"10",X"FB",X"18",X"B9",X"CD",X"BA",X"38",X"21",X"20",X"80",X"36",X"F3",
		X"54",X"5D",X"13",X"01",X"BF",X"03",X"ED",X"B0",X"21",X"8D",X"3E",X"06",X"0A",X"C5",X"5E",X"23",
		X"56",X"23",X"46",X"23",X"4E",X"23",X"7E",X"23",X"EB",X"CD",X"23",X"3A",X"EB",X"C1",X"10",X"ED",
		X"C3",X"A1",X"39",X"21",X"20",X"84",X"36",X"0C",X"54",X"5D",X"13",X"01",X"BF",X"03",X"ED",X"B0",
		X"C3",X"A1",X"39",X"C5",X"E5",X"77",X"23",X"10",X"FC",X"E1",X"0E",X"20",X"09",X"C1",X"0D",X"20",
		X"F2",X"C9",X"CD",X"AD",X"38",X"21",X"20",X"80",X"0E",X"1E",X"06",X"0F",X"C5",X"06",X"00",X"36",
		X"94",X"54",X"5D",X"23",X"36",X"93",X"23",X"EB",X"ED",X"B0",X"EB",X"0E",X"1E",X"36",X"96",X"54",
		X"5D",X"23",X"36",X"95",X"23",X"EB",X"ED",X"B0",X"EB",X"C1",X"10",X"E0",X"3A",X"00",X"D0",X"CB",
		X"4F",X"20",X"F9",X"C3",X"CD",X"35",X"08",X"84",X"80",X"52",X"41",X"4D",X"00",X"00",X"00",X"4F",
		X"4B",X"00",X"10",X"84",X"80",X"52",X"41",X"4D",X"00",X"00",X"00",X"4E",X"47",X"00",X"00",X"5D",
		X"00",X"00",X"00",X"00",X"5D",X"00",X"52",X"4F",X"4D",X"00",X"00",X"00",X"4F",X"4B",X"52",X"4F",
		X"4D",X"00",X"00",X"00",X"4E",X"47",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"36",X"21",X"37",
		X"AD",X"37",X"66",X"39",X"96",X"39",X"32",X"3A",X"B0",X"3A",X"B8",X"3A",X"03",X"00",X"03",X"04",
		X"00",X"04",X"08",X"0C",X"10",X"1B",X"26",X"31",X"01",X"73",X"81",X"35",X"01",X"73",X"81",X"33",
		X"01",X"73",X"81",X"32",X"01",X"73",X"81",X"31",X"08",X"ED",X"81",X"31",X"30",X"00",X"33",X"30",
		X"00",X"35",X"30",X"08",X"ED",X"81",X"32",X"30",X"00",X"34",X"30",X"00",X"36",X"30",X"08",X"ED",
		X"81",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"30",X"08",X"ED",X"81",X"00",X"00",X"00",X"00",
		X"00",X"00",X"4E",X"4F",X"FA",X"3A",X"FC",X"3A",X"01",X"00",X"00",X"0A",X"07",X"B1",X"82",X"54",
		X"41",X"42",X"4C",X"45",X"00",X"00",X"07",X"B1",X"82",X"55",X"50",X"52",X"49",X"47",X"48",X"54",
		X"16",X"84",X"80",X"44",X"49",X"50",X"00",X"53",X"57",X"00",X"31",X"00",X"32",X"00",X"33",X"00",
		X"34",X"00",X"35",X"00",X"36",X"00",X"37",X"00",X"38",X"03",X"C6",X"80",X"53",X"57",X"31",X"03",
		X"06",X"81",X"53",X"57",X"32",X"0B",X"64",X"81",X"50",X"41",X"54",X"52",X"4F",X"4C",X"00",X"43",
		X"41",X"52",X"53",X"0D",X"A4",X"81",X"45",X"58",X"54",X"45",X"4E",X"44",X"00",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"08",X"F6",X"81",X"54",X"48",X"4F",X"55",X"53",X"41",X"4E",X"44",X"09",X"24",
		X"82",X"43",X"4F",X"49",X"4E",X"00",X"4D",X"4F",X"44",X"45",X"09",X"A4",X"82",X"42",X"4F",X"44",
		X"59",X"00",X"54",X"59",X"50",X"45",X"00",X"01",X"2E",X"82",X"00",X"1A",X"64",X"82",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"9F",X"3B",X"AF",X"3B",X"00",
		X"10",X"20",X"30",X"40",X"50",X"60",X"60",X"70",X"80",X"90",X"A0",X"B0",X"60",X"60",X"C0",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"32",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"33",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"34",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"35",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"36",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",X"59",X"00",X"0D",
		X"31",X"82",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"32",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"33",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"34",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"35",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"36",X"50",X"4C",X"41",X"59",X"53",X"0D",
		X"31",X"82",X"00",X"46",X"52",X"45",X"45",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"2E",X"82",X"41",X"0B",X"64",X"82",X"43",X"4F",X"49",X"4E",X"00",X"4D",X"4F",X"44",X"45",X"00",
		X"42",X"00",X"03",X"00",X"03",X"04",X"9A",X"3C",X"A2",X"3C",X"00",X"10",X"20",X"30",X"40",X"50",
		X"60",X"70",X"0D",X"31",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"31",X"50",X"4C",X"41",
		X"59",X"00",X"0D",X"31",X"82",X"32",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",
		X"59",X"00",X"0D",X"31",X"82",X"33",X"43",X"4F",X"49",X"4E",X"53",X"00",X"31",X"50",X"4C",X"41",
		X"59",X"00",X"0D",X"31",X"82",X"00",X"46",X"52",X"45",X"45",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"32",X"50",X"4C",X"41",
		X"59",X"53",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"33",X"50",X"4C",X"41",
		X"59",X"53",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"35",X"50",X"4C",X"41",
		X"59",X"53",X"0D",X"71",X"82",X"31",X"43",X"4F",X"49",X"4E",X"00",X"00",X"36",X"50",X"4C",X"41",
		X"59",X"53",X"0F",X"8B",X"80",X"31",X"00",X"32",X"00",X"33",X"00",X"34",X"00",X"35",X"00",X"36",
		X"00",X"37",X"00",X"38",X"04",X"C4",X"80",X"4B",X"45",X"59",X"30",X"04",X"04",X"81",X"4B",X"45",
		X"59",X"31",X"04",X"44",X"81",X"4B",X"45",X"59",X"32",X"06",X"84",X"81",X"54",X"49",X"4D",X"49",
		X"4E",X"47",X"00",X"0E",X"01",X"00",X"00",X"00",X"01",X"10",X"11",X"12",X"13",X"14",X"16",X"17",
		X"18",X"1B",X"1C",X"1D",X"1E",X"1F",X"00",X"00",X"0B",X"27",X"80",X"53",X"00",X"4F",X"00",X"55",
		X"00",X"4E",X"00",X"44",X"00",X"53",X"0E",X"44",X"81",X"30",X"37",X"00",X"53",X"50",X"41",X"43",
		X"45",X"00",X"50",X"4C",X"41",X"4E",X"54",X"0D",X"64",X"81",X"30",X"38",X"00",X"55",X"46",X"4F",
		X"00",X"46",X"4C",X"59",X"49",X"4E",X"47",X"0C",X"84",X"80",X"30",X"31",X"00",X"45",X"58",X"50",
		X"4C",X"4F",X"53",X"49",X"4F",X"4E",X"0E",X"E4",X"80",X"30",X"34",X"00",X"43",X"41",X"52",X"00",
		X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"10",X"C4",X"80",X"30",X"33",X"00",X"55",X"46",X"4F",
		X"00",X"45",X"58",X"50",X"4C",X"4F",X"53",X"49",X"4F",X"4E",X"10",X"A4",X"80",X"30",X"32",X"00",
		X"50",X"4F",X"49",X"4E",X"54",X"00",X"50",X"41",X"53",X"53",X"41",X"47",X"45",X"07",X"04",X"81",
		X"30",X"35",X"00",X"43",X"4F",X"49",X"4E",X"0B",X"24",X"81",X"30",X"36",X"00",X"43",X"41",X"52",
		X"00",X"4A",X"55",X"4D",X"50",X"14",X"84",X"81",X"30",X"39",X"00",X"42",X"41",X"43",X"4B",X"00",
		X"47",X"52",X"4F",X"55",X"4E",X"44",X"00",X"4D",X"55",X"53",X"49",X"43",X"0F",X"A4",X"81",X"31",
		X"30",X"00",X"45",X"4E",X"44",X"49",X"4E",X"47",X"00",X"4D",X"55",X"53",X"49",X"43",X"10",X"C4",
		X"81",X"31",X"31",X"00",X"4F",X"50",X"45",X"4E",X"49",X"4E",X"47",X"00",X"4D",X"55",X"53",X"49",
		X"43",X"0F",X"E4",X"81",X"31",X"32",X"00",X"53",X"54",X"45",X"50",X"00",X"50",X"41",X"53",X"53",
		X"41",X"47",X"45",X"11",X"04",X"82",X"31",X"33",X"00",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",
		X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"10",X"24",X"82",X"31",X"34",X"00",X"43",X"41",X"52",
		X"00",X"45",X"58",X"50",X"4C",X"4F",X"53",X"49",X"4F",X"4E",X"00",X"00",X"00",X"A8",X"01",X"38",
		X"60",X"A8",X"41",X"38",X"98",X"90",X"81",X"38",X"60",X"90",X"C1",X"38",X"98",X"68",X"01",X"38",
		X"60",X"68",X"41",X"38",X"98",X"50",X"81",X"38",X"60",X"50",X"C1",X"38",X"98",X"20",X"84",X"20",
		X"07",X"00",X"00",X"87",X"20",X"07",X"08",X"00",X"85",X"20",X"08",X"02",X"00",X"86",X"05",X"08",
		X"05",X"05",X"86",X"04",X"08",X"0C",X"09",X"86",X"05",X"08",X"06",X"0E",X"86",X"04",X"08",X"04",
		X"12",X"86",X"05",X"08",X"03",X"17",X"86",X"04",X"08",X"00",X"1B",X"86",X"05",X"08",X"08",X"0E",
		X"84",X"80",X"30",X"31",X"00",X"00",X"44",X"49",X"50",X"00",X"53",X"57",X"49",X"54",X"43",X"48",
		X"0C",X"C4",X"80",X"30",X"32",X"00",X"00",X"49",X"3F",X"4F",X"00",X"50",X"4F",X"52",X"54",X"0A",
		X"04",X"81",X"30",X"33",X"00",X"00",X"53",X"4F",X"55",X"4E",X"44",X"53",X"0D",X"44",X"81",X"30",
		X"34",X"00",X"00",X"43",X"48",X"41",X"52",X"41",X"43",X"54",X"45",X"52",X"09",X"84",X"81",X"30",
		X"35",X"00",X"00",X"43",X"4F",X"4C",X"4F",X"52",X"0F",X"C4",X"81",X"30",X"36",X"00",X"00",X"42",
		X"45",X"41",X"4D",X"00",X"41",X"44",X"4A",X"55",X"53",X"54",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
