-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "193D1A0292A2AABBAEBA2AEA9A6BF50D844A4178BA4CD0FC21717FA329B9B7F3";
    attribute INIT_01 of inst : label is "210130DF1E20023FB2010DB67917D492927E6CC34D6A5350FB00EA2AAB1F7AF8";
    attribute INIT_02 of inst : label is "BDE1150552009416A045530284C0AA5028A1186C5534B3565ACB0186019A4C9B";
    attribute INIT_03 of inst : label is "2C0820101040011AC59C634331518A8C7473A39127F6F49DF0521F62B642CFA8";
    attribute INIT_04 of inst : label is "20BD9F4BF1A4C30C96D110432494092401040924000041000986192DA2208649";
    attribute INIT_05 of inst : label is "2101161FFBB8CAC1E5E135DA64D4449A9B06CB0F616C3FDE7D6DBB4A37E13744";
    attribute INIT_06 of inst : label is "2490208040410086E202D19B9412A8E85A72297E3684542E6CC1021438E2494B";
    attribute INIT_07 of inst : label is "9A0E619BE577CCC0820924802082492012480080820101040202082492008209";
    attribute INIT_08 of inst : label is "659EDC60AC2305140892E87111149213D6021414004400057695959594D76E3B";
    attribute INIT_09 of inst : label is "363091811188A28121DD214965B67D89202E252351BC8A0BA34993C8502C4A5D";
    attribute INIT_0A of inst : label is "94964CF5830DB364F649332D8806633018109662A2C93693E904F9CB93637B1B";
    attribute INIT_0B of inst : label is "32CEB30C80AF6ED6AB76B4F59BF6B75FB5A7AEDBB5AADDAD3D66FDADD7ED69EB";
    attribute INIT_0C of inst : label is "A6B624B0A26D437EE1BBDA1088569484961049286FC62632202C2901E800FAEA";
    attribute INIT_0D of inst : label is "DA86FF81B621BF96C377B42120B4A424B0E249437FE18D261B7D4F0DDC98C486";
    attribute INIT_0E of inst : label is "1760489A3D5421414466DD951532000219390EDF33A7B332B332802F5B125844";
    attribute INIT_0F of inst : label is "7FF803EBEABFEF7BE5836D36D37D77D76E6F2FAF2CAC02DCFB6DB6DA4ECDC897";
    attribute INIT_10 of inst : label is "A4E8C49286E6A661BCEE8CA380CEEC63CC718BAAAF2A6F26D76B0924B9CA2E19";
    attribute INIT_11 of inst : label is "9B89B50DBDCCC3F4992D18D271A7D449286D6A661F36E8C4DBA9B6E661A54D37";
    attribute INIT_12 of inst : label is "2373DC3C14494F4677755552AA9C0001FFFE0000FE9D2EB70BDE6DDAD18DBEA6";
    attribute INIT_13 of inst : label is "27FBB8C0B2BAB669D631D00E54846389B2AAEE4EEE01E04F0D0F0D0B090B090B";
    attribute INIT_14 of inst : label is "9F7E3EFC7DF8FBF1B7E36FC32A282FDF1FBE3F7C7EF8DDF1BBE40714572B88F6";
    attribute INIT_15 of inst : label is "8330660AA4A311102040811217805B6543AA36F739D868A6AC312D62A00CD19B";
    attribute INIT_16 of inst : label is "8A00005E05A398CC66902A40ACE61AB1CE64722294A3234414A55B6D248CCC19";
    attribute INIT_17 of inst : label is "6E26599B899766E26599B89975831F495754D4473D663D763D663D7364417C11";
    attribute INIT_18 of inst : label is "D93030BA418D6B044A028592A76432C10680A1A724975102A32635464C5C113F";
    attribute INIT_19 of inst : label is "36A4BB223B4BBD92B374D84FEEAA318F989DFB1761BB9264A2945B676EE8A516";
    attribute INIT_1A of inst : label is "9624962494490D53BBBA22227274D34D34B51B9BB92486EC6085A8282BDEDD11";
    attribute INIT_1B of inst : label is "DD973B11670A4AAA3263B8C3772490DDB31BB16F0A4AAA325B271DD3D8EBC824";
    attribute INIT_1C of inst : label is "B490DD973B316E0A0AAA3263B8C3772490DD931B91660A0AAA326338C377B490";
    attribute INIT_1D of inst : label is "8B4DB0431C908A538943F47C0203F0C60064C005FFFFFBEED5294B8EA3F8C377";
    attribute INIT_1E of inst : label is "BC20444194F3C29BA28D7884188488C49103108B6C4240B6C1C7243303881111";
    attribute INIT_1F of inst : label is "C2EA7E8C0A14A523FDB89B0DBB9009E339662013847AEE40278CE598804E11EB";
    attribute INIT_20 of inst : label is "90E91A0617742B01B2E0A6089DD2EDFD14C7BB68872FCC2AAA44F9FA7FCCF6C9";
    attribute INIT_21 of inst : label is "0AD3D1091E8DD34900103CB6A261427CA794EF24E04C2784BB498DD152E3A8E8";
    attribute INIT_22 of inst : label is "48971A4A829D6215A3744A0A0C42B468A8E89C38D68E886BA4DA3A258D146243";
    attribute INIT_23 of inst : label is "9921D1DB0D83E29E49D908214BAFFCC1FFFFFC3FFFFF0C01999E05E9934E9C4C";
    attribute INIT_24 of inst : label is "C3AE9193106FC74ADA9F73A97B5ED05094C4E80E72D6787B37E89C4FF7327324";
    attribute INIT_25 of inst : label is "97430F624BA1872125D2C30281A86A59F7B1497BB2125D0C358B7DDD6FB3A36E";
    attribute INIT_26 of inst : label is "BC90B288E228B17A64AE1C6EA2F9964924BD2C33165872125D0CBD892E961C84";
    attribute INIT_27 of inst : label is "995D92C9AFE7EE4B279DD9D2E9FB7A599CFCECE4B3E64B25ADC74A8B0B772B2D";
    attribute INIT_28 of inst : label is "C901F7974BA74BA35D92C992C8D674BA74BA75D92C992C95674BBE066CCF4B33";
    attribute INIT_29 of inst : label is "B22C27D3B9E81FF6B8E7EDDFF870C63DBCF8D73E3FF5203CD7B9FCF13259FE62";
    attribute INIT_2A of inst : label is "CD34D86432E0B48FBDB556D67EE11EF2BFC79DFF40C1A1081D3CCFB5624F9505";
    attribute INIT_2B of inst : label is "A4794679E7AAB4401F00C4A1F6D7FF7F032742EA7E01446294D80550404A5451";
    attribute INIT_2C of inst : label is "4CEC11A67508D33A6CE24DBDD85C77425B3F3E6AFD3F865F7A68AEDE9A37A102";
    attribute INIT_2D of inst : label is "A29A483050BDA8F6EE05B6B800007FFB603A9CCDD33B0C9E0106B155CEC533B5";
    attribute INIT_2E of inst : label is "7F8FFBBF0A5D362F9ADD2E3BF686E359E648D6C7BF5971A7FCF5D33B0EA2A2A2";
    attribute INIT_2F of inst : label is "F43D443ECCCE96B5EFFF3F5D4FD75375D4FD753EB53FFC850FA58576EEEEEEEB";
    attribute INIT_30 of inst : label is "0040000000002400000000000000000212400000600208000004024000000000";
    attribute INIT_31 of inst : label is "FB597D9E7287EAE9E6DBBFB40ECC912700000000001240040000000124A00000";
    attribute INIT_32 of inst : label is "1DA91D0018105CEC987BEFE9C7BCEC987B007FFF7FDD23C612FB0CB27E8E00F3";
    attribute INIT_33 of inst : label is "41F9FDFFD114662E62C444019F8BF1500C22E7A8001F188B89414787A2FAB333";
    attribute INIT_34 of inst : label is "800FB0DF0004000200424800038C70400000008048000000001C550467F2AF15";
    attribute INIT_35 of inst : label is "88A2222222088882208804000200024800830030002494038FF1C80001800004";
    attribute INIT_36 of inst : label is "DDF5D400023800007DF55DFDFDDDDDA23DD77772777DDF727775DC222228888D";
    attribute INIT_37 of inst : label is "0F6550A0000002177028E9388E90A61CA5D4F1F1C400F4E2F991C2ABDCD20D7D";
    attribute INIT_38 of inst : label is "751D4741D0761D07C7FEC1FEBBFE55C3F6AE5C1F6345C1F63059987079B607B0";
    attribute INIT_39 of inst : label is "A7569DF6EFDB81CCCE4A77D3B53D1A9C06193D507672AAE4E551D9E029F2F9D4";
    attribute INIT_3A of inst : label is "A1958850FFF50078F001FEF17C3DDFBF800F00001E3FBFD50FFA87F6A5FBF2EF";
    attribute INIT_3B of inst : label is "1294249FF11FE0B0BA01F28E1A432452442C00000C484C4CD041FFFB1C471F03";
    attribute INIT_3C of inst : label is "CCFF79D3FFFFFF25804631DEC47CAF2AD0B050023FD50DAFFFFFFDA494A5014A";
    attribute INIT_3D of inst : label is "7406E6701A9D806B7E01644E77860B6899B3E205A44E9E44F5DEA6B74897A3FF";
    attribute INIT_3E of inst : label is "DB0FAF9B7DB2009900893449BDC0CE4266D7B951515101BE2A2A6CD4F90FFC6A";
    attribute INIT_3F of inst : label is "D5749BB762CC99733CEF5A675CCF3BC6939243930F3259993201F7A4D50BA42D";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "3267A0FD2FD77DE4DA6DB69A7DF7BBD6027D68278718A22F7D69911BD5DF5F8F";
    attribute INIT_01 of inst : label is "63AD7C2502D09340216CB26425A100240C8082FBAED93526576417C7452AE30B";
    attribute INIT_02 of inst : label is "5B5FEB53A9CF9FBCDAFDA437D53BFF73FFC577A9270E24801080E830AABF5E23";
    attribute INIT_03 of inst : label is "40530648820493C0CC18C25926223113888C449B3774EBD697F7B104473EBFEE";
    attribute INIT_04 of inst : label is "5B6178B482221A202088A60A08225041882050418922081244344041114C1410";
    attribute INIT_05 of inst : label is "7CD8C979144300061F4E4D24A9A99D3562F192D45E8B434986192685C908C5BF";
    attribute INIT_06 of inst : label is "00014C1922983247097FE231BB7F998EA5E4D749EDBE9F6DB0C2F4CBE51984B4";
    attribute INIT_07 of inst : label is "6C10CEE21E09F34410400011041000048001324530648A60C910410000441040";
    attribute INIT_08 of inst : label is "DB2891D2CF8F24AFA8B2482ACA414DF8F8000155112708B04022828280228180";
    attribute INIT_09 of inst : label is "4887035B415C95F51589BB1925B2C954DB755ADC4132D3EA0253E9BEDA8BAD06";
    attribute INIT_0A of inst : label is "DB99E55D75D0004AA4928CD979F0C99DB5B225AD2DB6D26D21A9432064B0A735";
    attribute INIT_0B of inst : label is "6C799641FF42BD4BF5CA4D596D5ACDEAD66AC9AB52ED5293564B76B3FBB59AB2";
    attribute INIT_0C of inst : label is "5949CB063593B090D84027396569293B21C29272020C8CA56D72F36A8EAE40B8";
    attribute INIT_0D of inst : label is "6F6120F2DBD84C7B3080DC62CA5B5BD90E34B79010DED2DC80C3B6402371892B";
    attribute INIT_0E of inst : label is "8816AB4DA0DE0C5D31D8B56662589FEDB625D320B54846EECAC52A81ADE5830B";
    attribute INIT_0F of inst : label is "83100115C1C09C86958124904134D145A23E5E5ED504A488C6DB6DB6DDBB004E";
    attribute INIT_10 of inst : label is "C997892520340A0D10B50B42509333302604C2DEFFFCB24B6886404126296983";
    attribute INIT_11 of inst : label is "C116DAC210943A4B76D2D12D965D0896D20084A0D249B38B2492680A1D71B240";
    attribute INIT_12 of inst : label is "580532D22FC280AA0CFFFFFDFF92000001FFFE00213640E49F25B76D6516D2DB";
    attribute INIT_13 of inst : label is "0A4ECC7F491568F669C62FF1A8AA9C7267C51114196F093A78787A7A78787A7A";
    attribute INIT_14 of inst : label is "51ADE1D946B787655ADE9D90F65F696AF274A5ABC9D2B6AF674EA12F8581624B";
    attribute INIT_15 of inst : label is "1666CCC3B23022224599166A60B58A0C9ACD187FEB128B4CCB664A2DAFA9012E";
    attribute INIT_16 of inst : label is "3CC9C8B79E4CE330B84E691BA514A5617E97D49B0BB5C5B9D85DE4B2F9108891";
    attribute INIT_17 of inst : label is "9188D2A4E274A9188D6A4E27582A40E7C0D9A412D24AD64AD25AD65C5726DE26";
    attribute INIT_18 of inst : label is "72D290459BDEF724CD6D6927CE49F9CB355B5AD7386ABEF81CC8B03991761A7A";
    attribute INIT_19 of inst : label is "08D36CDAC5BE59612CC8232800DAC82225C444B8C800248B2724E4CFE809C939";
    attribute INIT_1A of inst : label is "2D2B3D2B3E567EF84C4C4C4C04C96CB25B5D6480024B611060EE7D73F17E0686";
    attribute INIT_1B of inst : label is "0043124BB3DDDD01CC8A441000496C220312EB9BDCDC01CC9A4C4B24B6B15F2B";
    attribute INIT_1C of inst : label is "DB24004732CBB2DD9D01CC8AC41000D96C2247324B92DC9C01CC8ACC30884B24";
    attribute INIT_1D of inst : label is "34280410532C14D9B6670F83FDFC0F3DFF9B3FFA0000F209BFD0B554500C3088";
    attribute INIT_1E of inst : label is "56BD37BD7B07052E26BC933583445512C818363541105B141114CB02AEB36693";
    attribute INIT_1F of inst : label is "03D00009057BFEFFC3A67AE7ACCDF3BDE3498BEF7BCEB137CE739D622FBCE71A";
    attribute INIT_20 of inst : label is "3AB68F4DE59ED46A4C0F58E6628D121AEB3B44D4E800012AAAD50FFAFE602952";
    attribute INIT_21 of inst : label is "5326645719126DB6332B8069C83CB4995B7B6A4916E3DB3B6D9232652D411F34";
    attribute INIT_22 of inst : label is "E365A59161E290E6489915F47E89E4499111023935511196C91544566AAE90B0";
    attribute INIT_23 of inst : label is "0809C4AE2F1FEF15547EE5A5F41000FFFFFC003FFFFCFC0181FCE70840800106";
    attribute INIT_24 of inst : label is "339E3880DE3F0C21804421440005090A00294C018C610524D9BB6D024C102101";
    attribute INIT_25 of inst : label is "30B44094B8CE604EC82F10FD6AF795A4481402C544EC82D10A585B430B605848";
    attribute INIT_26 of inst : label is "FDC2F57DFDF925FD4F51EF05755429965922F106E18604EC82F106F2C329836B";
    attribute INIT_27 of inst : label is "91766D37AA09D1B4DC95F625130F84A244BF910B4498B4CAB13608773F2F575C";
    attribute INIT_28 of inst : label is "36C0D06994C994CC766D366D370D894489448722D162D178C994C89A10D1945C";
    attribute INIT_29 of inst : label is "4C4249A463B34A9B274C12004B0C395261C764CF551A52A72863D78EC5A3EC15";
    attribute INIT_2A of inst : label is "34D34B2926A4C777E592DA4532C7EFB143EFFFDE36EDF7FDAC03E80A9C9C6252";
    attribute INIT_2B of inst : label is "F2FBF40102FFC6FCBE3D2F3E34D40E5C4CCC36F139DD2A89CDF8044401232DDB";
    attribute INIT_2C of inst : label is "A2239B19128D88890825702454E614721978001F15FF96FBC8FEEE5A34D71397";
    attribute INIT_2D of inst : label is "4CEAAD4CA76CCCB3E8CE42F00000775C244F660B5C3159AC580BCBEB203AC88A";
    attribute INIT_2E of inst : label is "B7A2F01F1CF2D27565965455215CBCD2E0540A4EFEB25E0381F35C315ACC44CC";
    attribute INIT_2F of inst : label is "CFD0DB01A510400053FE8D27B149EC527B349ECDEEC002C99636499AFAFAFEFF";
    attribute INIT_30 of inst : label is "413B6080417B65ED824905ED824905ED8009DF20D04BBE416093B6DEEFFEFFEC";
    attribute INIT_31 of inst : label is "86961968584E1494C02A401003266C4C0D824105ED800BDB27FE49DE183B6080";
    attribute INIT_32 of inst : label is "40883FA4C81BC1A153003A357043B35700007FFDA44686BC0182E02DA1490044";
    attribute INIT_33 of inst : label is "0A061201E14209D19D5051EA60741441021D185000008274664450781D052121";
    attribute INIT_34 of inst : label is "BDB86BB0BDB05D73BDB4933BEE7A0B76EC2E1A76DBDDFFDFFD9E502A184D5794";
    attribute INIT_35 of inst : label is "DDFD7D7D7D5DF5FD7F70B44831BDB4037B76FFED3BCB276E7808276E190C2F6D";
    attribute INIT_36 of inst : label is "0A82A88882922222555FF7E055555F57D5FD7FFFD7D5F5557FFF5FD7D7D5F775";
    attribute INIT_37 of inst : label is "6E0996E0000003138166A3406F8924DC456C19720CFCAD06E0A9C06BBC95708A";
    attribute INIT_38 of inst : label is "7ADE77ADC372DCB737FE69F5218A99C1D349DC1C3459C1D340CA0F70F0E86340";
    attribute INIT_39 of inst : label is "578B56CAB5AB8DCA6E137993AFBB97DC00073C34B270636CE0C2C9C819F189E7";
    attribute INIT_3A of inst : label is "B722D424910AAF85156A2115C00004043F10F8BE21E23FAB6FDEB5F42D7516F7";
    attribute INIT_3B of inst : label is "4FBE8040172F2F9F9202E8C3736688A04C0C444144404F44D861FFAE10A10C9E";
    attribute INIT_3C of inst : label is "C00068D03FFFFE88401085319A18B6349D0B9372D31D953FFFFFFD8127EFAFDF";
    attribute INIT_3D of inst : label is "8C1B69D865A761B4B1C0B7994A6B04BF76ED3D82DF9B7A005F991925AB023C1D";
    attribute INIT_3E of inst : label is "327F54BD0FD7FEF400525A92C001613000781C04040300006EE4932910D3FD94";
    attribute INIT_3F of inst : label is "04DF0674B51B26C51B890859B166F2421C65902E606CA8320D000449E5D64913";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "38714DCC6724B2CB2CB2C92CA2884CC8B8944C4A28A208111E28363680B66868";
    attribute INIT_01 of inst : label is "522A5F02E0108302D3B58DBF5985B508A92B84924954AE3A95C613266652A13E";
    attribute INIT_02 of inst : label is "DAD5ED7A230C552694E58C73C307BE1FBE21571DE21880901282B73E02FFFF48";
    attribute INIT_03 of inst : label is "DA24D134492248004C48C74603331998ECC766385C09868329898A28863AEFEF";
    attribute INIT_04 of inst : label is "99A5D57F5A21B49A6D256D26926D26934492349344912489236934DA4ADA4D24";
    attribute INIT_05 of inst : label is "31D8B8CC275A01E8B57335CE67B304F63DB4CD39A33462FFFBF5BCC91560F723";
    attribute INIT_06 of inst : label is "92489344D12689A819A491619DB49DC22FB41DF3AD36592B9CA0EE8B8A3D86CB";
    attribute INIT_07 of inst : label is "749A7C53347D6B424924924892492492492489A24D13449A2689249249224924";
    attribute INIT_08 of inst : label is "3ED6DBB287CA08263992F82CD8E54925B8800001C99681B910A5A5A5A56AC1C3";
    attribute INIT_09 of inst : label is "05D3816DE36504C7B05F99C96C92494449BD98C6B3E4EB2F47CF60265DDE2DFB";
    attribute INIT_0A of inst : label is "A34DB0E1D6189972525B99C043CB9DDED6DF2AE928E3893C159D1835DA608C13";
    attribute INIT_0B of inst : label is "BA8E23A50C4EC5CF060E6CE59EBEFA74F7672C70F74387BB3961839A0C1CD9CB";
    attribute INIT_0C of inst : label is "6474661B4E4CC32B21999BBD918C8E8EC269CD186566373929634D4B272BC2EB";
    attribute INIT_0D of inst : label is "D1C75513B471D18C63BB377BA26474641B4F68E3AB231DA71D58C98ECCDDEECC";
    attribute INIT_0E of inst : label is "C2BB286A89580E4555456982339CA9B4D7B8C482636DD712E3918AF23A3A099E";
    attribute INIT_0F of inst : label is "96C8E0DB09616354E981F7DF7DE79E798A191919179B3A12FFFFFFFFB12DB696";
    attribute INIT_10 of inst : label is "B4C98CD18651C7A641E55E0781E4E6C2D85B0B1AE4BA3DFDB263996DB89B1A0D";
    attribute INIT_11 of inst : label is "F71DA38E738F6C269D1D91DA0136B8ED1C739C7B6134CD8CD009B5C7A658DB7B";
    attribute INIT_12 of inst : label is "5CE3CD1326534366330AAAA82ABC00015555555454D998262B8269D1D31DA026";
    attribute INIT_13 of inst : label is "07B9982ECF9104B11CD9A2DC48E2C0C3DB17FB8C669A0990525252D250D050D0";
    attribute INIT_14 of inst : label is "BA76346C6CDDDBBBA76346C9F64CDD9D1B1A3736EEEDD9D1B1A6B3260E0783E6";
    attribute INIT_15 of inst : label is "E9D9B300B780CCCD1336688A823A2224EB912E914259C420600321312AFCE1D3";
    attribute INIT_16 of inst : label is "BE0C9D899F06B95DAE7449D1270647BF9EC26611DCB06ECC8EE5CA6DEECB674E";
    attribute INIT_17 of inst : label is "1C0E1DC7038771E0F1DC783C74FB8AB0B359E464387738773C773C7476722663";
    attribute INIT_18 of inst : label is "18A280D761084200607060D284344082141C1990187299B633A20E46665807A4";
    attribute INIT_19 of inst : label is "F8C4791A136B7583BA5FE32E76C221954BEAA17D619D98760F81F1670F43E07C";
    attribute INIT_1A of inst : label is "C84ECA4ED49D90AC6EE77FF73276924936667919D9B68674609F20F8BD2E1CDE";
    attribute INIT_1B of inst : label is "EC923B27C8BE2F72333390C33B36D0CED23B87C0BE2F633A139CC18C58C72C4E";
    attribute INIT_1C of inst : label is "34D0CE923B27E9BF6E72333398E3B33498ECB23B27E9BF6E633A2390C33B3698";
    attribute INIT_1D of inst : label is "C0A8104516D186508843FAFEF6D3F9E360ECCAF5FFFFFC276AE2D8CE67D8E3B3";
    attribute INIT_1E of inst : label is "171E3BDEE747099CA88FF445544567C0901A17404444544442C5B40ACFC48894";
    attribute INIT_1F of inst : label is "4358214E0262388E7DB8D3ADB910CDE62D722193CC52C4632798A588C66F314B";
    attribute INIT_20 of inst : label is "DAEC93576622C831380775B21938DED288E86646648C019154DDEF56D56CADDB";
    attribute INIT_21 of inst : label is "1B8ED239099F9245545551239C79C6C0E05C0F36FB4AE01C56DB77D331040E64";
    attribute INIT_22 of inst : label is "6B82324B90F8CC7719F48E2AAE3DA0C099DDF23181999DC56D9777630334CA64";
    attribute INIT_23 of inst : label is "584C4E1E2F17E84A58F8C0A103A00F01FFFC03FFFFFCFC001E1C761C2021038E";
    attribute INIT_24 of inst : label is "73163DA89A17005214E15AC84211891607BDEC0310C40E8C0668851466B8AB41";
    attribute INIT_25 of inst : label is "9361B346693099A3B0904CDEF718C5FFB6E44496DA3B0934CD917FCE2FF9D97E";
    attribute INIT_26 of inst : label is "7DA77631FD9835FC6F1599253165DB6924C9245AB3681A3B09244D1D0683668C";
    attribute INIT_27 of inst : label is "181CD1ECBB350347B21C9CD1EC1C1A3D90E6E6B67A63673405914A4713AF674C";
    attribute INIT_28 of inst : label is "1745E3CB67A367A41CD1ECD1EC07347B347B45CD9E8D9E817367A6060C036732";
    attribute INIT_29 of inst : label is "72606D36ABC1F966D4F14CCFD370AE76AED99395E2A362B5DAABE2739B3DE3DE";
    attribute INIT_2A of inst : label is "326A2B3D94A6C19F814A41110A24C0CF01EBCE2A30080C211809F0E048DC1323";
    attribute INIT_2B of inst : label is "C4FB9D44615540F93E3BB9BC2DB58A576E13321B429D63DD69000504043321D8";
    attribute INIT_2C of inst : label is "F7431DF3AA2EFDD0314670B49F68A67208599B3791FF16F580F443203E416CA7";
    attribute INIT_2D of inst : label is "E6BAF4E8F7F8CDE3EA8B74FAAAAAD7FFA477FDECC6085EBD12A5499F74379D09";
    attribute INIT_2E of inst : label is "DFDBFB9F16FFF45DB7FFFB6EFFDBFF9B8659DECBFEFFFF2035F4C6085A6666EE";
    attribute INIT_2F of inst : label is "89155602C84485211BFEE7FBF9FEFEFFBF9FEFEF7FE002F4E7B771DFAAFFABBA";
    attribute INIT_30 of inst : label is "BEC4DF7FBEC4DB137DB6FB137DB6FB117FF622DF6FB44DBEDF6C4DB110010010";
    attribute INIT_31 of inst : label is "FA5CDDCB7006E4E7879A322406C999A9137DBCFB137F7622D801B623E7C45F7F";
    attribute INIT_32 of inst : label is "083001203B6C86BE5D194BC591D4BC591D007FFCCA892AEE0B4B8BB9EE6E0016";
    attribute INIT_33 of inst : label is "B5FBEFFFFD69362EEA8F5A159F8BFC623162E7A800004D8B98C44007E2FAA121";
    attribute INIT_34 of inst : label is "6268B6D16268B6D3622FFEC45A6D1688B45A2D89B6220020021F96D16FBAAFE5";
    attribute INIT_35 of inst : label is "88802A802A8880A028036CB791626FEEC45B0036C47CF88A6814589A2914589B";
    attribute INIT_36 of inst : label is "8A0080A0A800A0A0F57D554200000A82AA0A8000280A02AAAAA80A0282A0AAA8";
    attribute INIT_37 of inst : label is "8A0E18A0000001164820E7240FF24255F15CD5F92000FC90E4E1C583D08A8280";
    attribute INIT_38 of inst : label is "5C1745E1585415058500C14A0964D5A017335A217555A007641A446801DCC2E4";
    attribute INIT_39 of inst : label is "D7B75E38FAA381E8AE657A4B9C3F8E1C011A3AC0A0758140EB0281E045D0F578";
    attribute INIT_3A of inst : label is "2D061C61000054020AB4010E45862040E1E00F43C00038002E2B970941CB40F1";
    attribute INIT_3B of inst : label is "9637206FE11F9B207604EC061242EC21444C054108484848FC48FF44B96E5B23";
    attribute INIT_3C of inst : label is "42705EB1FFFFFE2FC15AD7AD83D685B14C5CD59A3A800D0FFFFFFD2A458DC31B";
    attribute INIT_3D of inst : label is "F40C9F603A7D80E5EE41C74E75DC0F4E9D3AEE07A76E9440CA8D3B06885CBC15";
    attribute INIT_3E of inst : label is "AB314CBE383718B8004D20200000C77006F8808AA8040048C46724CBE0F3F065";
    attribute INIT_3F of inst : label is "149745B724E48CD315EB0A7334C5FAC29ADA40D1A9921A8819003307B0C5741C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "2B22CC3FF00800000000000000004ADBBE912440000000103602EE0A240820B0";
    attribute INIT_01 of inst : label is "3A0674104A101D42F3B1AD965AA4B508A9345904100686B604549F4E6640859A";
    attribute INIT_02 of inst : label is "DCB06E1BF586C57610FAF65A7595255D25650FDD8A1A841412807FDEA941A360";
    attribute INIT_03 of inst : label is "009244900000020A8BC4201A1111888C4462232A0A03572961A5A2A22E1ED7EA";
    attribute INIT_04 of inst : label is "192EF6F941E00041000000904900924800008248000000000000820000012092";
    attribute INIT_05 of inst : label is "1E775232448CBC97653366B606AD08D5B4D55148290526FBCDF4940F2FF073E3";
    attribute INIT_06 of inst : label is "00024912449224882924F1A0393CB5A23296997B927AAF2E4E72FF13E9F77938";
    attribute INIT_07 of inst : label is "0F95B98C48B2C440000000000000000000002489244912489200000000000000";
    attribute INIT_08 of inst : label is "B6D64EE2E699303A803248399B456DABDC008888E5CF01951AA5252525411B09";
    attribute INIT_09 of inst : label is "1E9980ED40C60750745B5B59249249C4692F3CFB70765157A0CD3B66CA862BFD";
    attribute INIT_0A of inst : label is "779FF0BEB318D92E5259DDA6E5F689C6DED21B618777887886BC9C65DB40DA1A";
    attribute INIT_0B of inst : label is "5CF735E48DA562BD8B15E8BEE3856E1C2B45F71C2B70E15A2FB8C15B060AD17D";
    attribute INIT_0C of inst : label is "6C76641B66ECC323A199DFBFB1ED8ECE8368DD986462A2968944204A868EFB73";
    attribute INIT_0D of inst : label is "D9864713766191CDC333BF7F636C76661B46ECC323231BB6195CD90CCEF5BDCD";
    attribute INIT_0E of inst : label is "13BB23CBAC4E261C3C7F6CE2AB7C0934DD14DC82722F93156971A3A63B33098D";
    attribute INIT_0F of inst : label is "BCF802C60B3553FCB883451451555554E40191919C81AE112924924926D24922";
    attribute INIT_10 of inst : label is "34CD8DD98642C52A55755755C17EEEEBDD7BADFB7DDFDBF7D32D4B6494DF7E09";
    attribute INIT_11 of inst : label is "BB1BB30CB58A54369D9991BB01B5D8DD9865AC42A1B4CD8DD80DAEC42AB8493B";
    attribute INIT_12 of inst : label is "CD428BB2BAC64624A2822222802A000067986798BC9D6852AAA369D9931BB036";
    attribute INIT_13 of inst : label is "0571703FD86FCB7AF3A25924F5FD2F2C8D66510945D85982C2C242C2C04040C0";
    attribute INIT_14 of inst : label is "6AD6D7AFAB5A54B4A96952D91C7555B56BEBD6D52D2A5A54B4A9F2BACACCB12C";
    attribute INIT_15 of inst : label is "D99D7F48C7A1CFCF9E2C58AD8B3620ACD15B3C08E60A26D656F3521DD55520A9";
    attribute INIT_16 of inst : label is "53ECBAEFE9EBD5EAF5B546D518C2EE9EBF5B2EDA975E3E47D4BABB4936AE777F";
    attribute INIT_17 of inst : label is "CDA68EF369A3ACDA68EF369A3E8953F6126CC849AB3BAB3AAB3BAB3A3EEBAFB5";
    attribute INIT_18 of inst : label is "FB1040927FF7BF38C66F6CD2E3344ECC2B9BDB9C2E3AFBBB2777C66FEFEE2B41";
    attribute INIT_19 of inst : label is "AD765794FE496EF8D7EEB12F7774F3C8B53336A6E9DD9EB594F29EEF8F653CA7";
    attribute INIT_1A of inst : label is "C984C984D70993FCA223B3333364926DA4743E1DD9F586642089E74FDDC998D4";
    attribute INIT_1B of inst : label is "ECB6B5E25952F6227669F1C333BCF8EE96B5725DD2D6327751ED4AB4AA5B5584";
    attribute INIT_1C of inst : label is "BEB0CC96B5E25952F7337F79F1C33BBEB8EC96B5F25DD2D7237E69F1C333BCB8";
    attribute INIT_1D of inst : label is "C884546134938498374305210B2C561C9F13350A0000F43648E8F98A7631C33B";
    attribute INIT_1E of inst : label is "6B2F1ADEA7E2E11085313E78B54ACDE40098136825608C0050CD2412CFE78AAE";
    attribute INIT_1F of inst : label is "411845250A52B4AF7D5FD5DDDFB8D967A9AF71B2CF535EC3659EA6BD86EB3D4D";
    attribute INIT_20 of inst : label is "E258DC42EAE3DDCED7BAB8C4CE07243F1E119364E70644AAAA0C95FE7FA4C5CB";
    attribute INIT_21 of inst : label is "35B4922FA08900054551410368117B50AA15413E3B68AA17DB6DA1931C4515C6";
    attribute INIT_22 of inst : label is "5EA25656BB78CC6F6C6483A2A3C9210308CC9160ACCCCD5DB6E2222551115660";
    attribute INIT_23 of inst : label is "D80834DA3D52F18A988E47CE2A88000000000000000000000002AF85402A0503";
    attribute INIT_24 of inst : label is "431C1D80BBE4434290C41AA842158DD38EBDB40EF7BD5F4A9C13584033B03B01";
    attribute INIT_25 of inst : label is "D2690766493483B3A098496B5AD6B6DB6DA654823A330D1694B3368866D113B4";
    attribute INIT_26 of inst : label is "3FA33E99EC81937D2546112731C68E49265D269B3A783A330D361D9984824ECC";
    attribute INIT_27 of inst : label is "0C8FD2FF19FE874BFA0A4FD2FFF43A5FF0527EF6BFFF6BFE40F358C23284C2C2";
    attribute INIT_28 of inst : label is "3F43EB8F4FEF4BECAFD3FFD2FF3BF4FFF4BFCEFDBFFDAFE2BF4BFED43D274B7E";
    attribute INIT_29 of inst : label is "6A3C2F97A97D51759AAD7CCAA130DF26ACD9D3B0F2F9783BFBA93173BA5FFF5E";
    attribute INIT_2A of inst : label is "A0EA0D3C5555A7FFD243E051BCCE61EF7E2A61FCB70E56B5D01D57BF7B9B51E1";
    attribute INIT_2B of inst : label is "5078AE640244505C1F9F983F0B2441407467B5FE73CEA888E4D0000110653A8A";
    attribute INIT_2C of inst : label is "F7666EB3BA575DDCA2C3FD998EA963FC287B8E26242FCC4C7C4570EF12F08082";
    attribute INIT_2D of inst : label is "A330E72A73D6BB501AB7F59AAAAAFD499474B97887B16D3F12A919DE74679D99";
    attribute INIT_2E of inst : label is "CFC9F9AFC669F4BADF496EBB95B76789EABD5695BDEBB3281888C7B16E2222AA";
    attribute INIT_2F of inst : label is "F93D5617CAE684215BFFFA4A5E929724A5C92973197FFD2E5DE72FFEAAFFFBE9";
    attribute INIT_30 of inst : label is "BE5D5F7FBE5D7D757DB6F9757DB6F9776DB2F2DF6FB1FDBE5F67F6DE30030030";
    attribute INIT_31 of inst : label is "BB6E74FE3A07E479E7D0FB240C899123157CBCF9756532EED805B2EAC31DDF7F";
    attribute INIT_32 of inst : label is "019C0984514CECFC4B39CEC4B3DCFC4B3D007FFE58AFA37E1A5DCE9FEE6700BB";
    attribute INIT_33 of inst : label is "A00DFDFFF680C1D33505A000607402DCC095185000003054650D280015052121";
    attribute INIT_34 of inst : label is "AEAFB2DF2EA3965F2EE4925C4BEC723FB7CBECFEDBC60060061F6A80B7F557DA";
    attribute INIT_35 of inst : label is "88802A802A88AA0A82AB23979F2EA4A25DDB00B65C4823BBEFF1CBABEF77CBAD";
    attribute INIT_36 of inst : label is "D55FFD77D817F55FAA22A0002AAAA028000000002AAAAAAA8002A0A8280A0000";
    attribute INIT_37 of inst : label is "2ACFFAA0000000122820AF140B80085515444160A4FCAC52F4A5C20B9167FFD7";
    attribute INIT_38 of inst : label is "5F1785C14050140505FEC570C9A09181C286181C250183C2180B006070830218";
    attribute INIT_39 of inst : label is "95085592A48B85D42E217B0B8CBB865C0500B900E17201C2E40385E001F2D17C";
    attribute INIT_3A of inst : label is "53061C600008040010200000024200000000000000002FC42BDA95F3857072AD";
    attribute INIT_3B of inst : label is "C73BA065010F056AA408F8861A43E4308C40480E04404444E468FF881EF21A5A";
    attribute INIT_3C of inst : label is "040837203FFFFFA100C6308CD3741D1F4DDCA394EED1E93FFFFFFC2A45CEEB9D";
    attribute INIT_3D of inst : label is "740DD770365D80DECE41DAC73FCE0EF5CF9FE6076AC78040B2C5B326E3D6590A";
    attribute INIT_3E of inst : label is "E9E6498A0723DF7800801400A706815032F42A0A222201505776FE8EB7DBE047";
    attribute INIT_3F of inst : label is "153B89ABE2DD9CF21DEA8F2F3C877AA3CF9241B32F76508B1101B7E698DF6604";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "237486209800000000000000000048987BB03300000000097AA808284600A205";
    attribute INIT_01 of inst : label is "42D5461A87515052E4C9280D942028750600040000112426755404C3700EA082";
    attribute INIT_02 of inst : label is "187603608C59E83550C82824921249124957BC9032D72EA1C4B8021000C16286";
    attribute INIT_03 of inst : label is "9324992649324D50296846280333199AEED7764690001122052122B760A53063";
    attribute INIT_04 of inst : label is "D6D8303209792492492649249249249264932492649924C9324924924C924924";
    attribute INIT_05 of inst : label is "FD820B20440001300718D860221A0443001330C018030349820360944180408A";
    attribute INIT_06 of inst : label is "924C92649924C93550490041A6CB1115A88556A05209C2C0088A94024559E480";
    attribute INIT_07 of inst : label is "4A727F20940013F24924924C924924924924C9324992649324C9249249324924";
    attribute INIT_08 of inst : label is "080DB1474908AA8999A400429288301000A8A0A073F2899A0D08080809128588";
    attribute INIT_09 of inst : label is "2101013283155133241213920024001696505210E342384246840824C701A802";
    attribute INIT_0A of inst : label is "4B0D87042699110956DB511003815003232C041D1C0A282200680182480092A4";
    attribute INIT_0B of inst : label is "05A16844098CD18D56AC7B04268C6AB563D8213063458B1EC109A31AAD58F608";
    attribute INIT_0C of inst : label is "4949420024928032801126332149292A400492500650D984E9D1974E24AB0616";
    attribute INIT_0D of inst : label is "250064524940190900224E764249494200249280328A924801D494008939D90A";
    attribute INIT_0E of inst : label is "400CA501B3860A28E3888073324076CB62049240E46F160048442AC0A4A10409";
    attribute INIT_0F of inst : label is "12300001101099401900820820924925A648585850006744D492492490092490";
    attribute INIT_10 of inst : label is "49200925006108C2F81AC1B0781191923246484C398D22D268D874DA07127106";
    attribute INIT_11 of inst : label is "04124A004213810922542324CE4820925002109C2849200926724108C040DB62";
    attribute INIT_12 of inst : label is "D4840062099E00A8C077D7D77F820001E1E1E1E0432254219E709225483249C9";
    attribute INIT_13 of inst : label is "08C88849506404EA515217A0210A8429C8D4AA91803E68B37173F173737173F1";
    attribute INIT_14 of inst : label is "79F1F1E1E3C3C7878F0F1E114413DC7CF878F0F1E1E3C3C7878A220990A2288A";
    attribute INIT_15 of inst : label is "0020040509402222448912210324000898454A5DF78201486342E2241AF36030";
    attribute INIT_16 of inst : label is "50BAEA9CA856351A8D49852614A085BD901B64D99B8576EECCDC26DBEDD80801";
    attribute INIT_17 of inst : label is "D96CC2365B308D96CC2765B308804093A88D8019440844084409440C0BAA72AB";
    attribute INIT_18 of inst : label is "A78220102D4350B2D7CE4E4DB593662CA3F392D8EB2826CC4000488000862261";
    attribute INIT_19 of inst : label is "543344D14890407C8549526156315208B1311E2798156F10C438879F41610C21";
    attribute INIT_1A of inst : label is "6C806C806D00D881777777762C9B6D9249402E0156D0414440485643152D22AA";
    attribute INIT_1B of inst : label is "08E080721D10E544000049002A4A400A8080721D10C555092050AC2A82156380";
    attribute INIT_1C of inst : label is "4A0828E080621990C555091049002A4A0008E080621990E554011049002A4A00";
    attribute INIT_1D of inst : label is "06030404000156385CB5F67EF4B3F3EDF364CFF5FFFFF49182A94913AC89002A";
    attribute INIT_1E of inst : label is "D3EF9B9EE700352316537112A103150920BCAD04110428001000000C68112249";
    attribute INIT_1F of inst : label is "43543301035AD6B5060D68F68C689110E618D12221CC31A24443986344A88730";
    attribute INIT_20 of inst : label is "6A36ED51808BB4614C8D50E6B01002026D3C0404E92100440019A5545520058B";
    attribute INIT_21 of inst : label is "B328669689986DB40011100A5025B902D84B02DA0CB2D85B0DA440662C501137";
    attribute INIT_22 of inst : label is "9B69A59978E69D665019A5AA20B048D09999E11939999990D266667673359500";
    attribute INIT_23 of inst : label is "4008A8B0F070116A189AC28427200000000000000000000000014D3F83BC1A04";
    attribute INIT_24 of inst : label is "41180C019B962810043010C318C28985933BC405AD6B13008825062000800801";
    attribute INIT_25 of inst : label is "510830942880084A9040040842108400000681C64DA104A0027FED89FDB13FEC";
    attribute INIT_26 of inst : label is "02630904B085380370D42608452478001044B04C20240DA10490425082506128";
    attribute INIT_27 of inst : label is "804620105592A8800B820620108444007C10310A0580A00B48724B30AA00B0B8";
    attribute INIT_28 of inst : label is "B6C04A288450805142211020114088440804142291028105088059184228808B";
    attribute INIT_29 of inst : label is "65372D13EB3161592301408A91000B42E8CC6494D29922056BEB50188C07EDBC";
    attribute INIT_2A of inst : label is "084880080C501C404040A860434E0E1EC18B290A256AAD6BA02154C12C482999";
    attribute INIT_2B of inst : label is "3304696684414705C04508326FB71B765208271585A88954204D100400000E46";
    attribute INIT_2C of inst : label is "0571C60AB1C10119C6C637B79CAB66342A5FAE3706802804081DD02205481298";
    attribute INIT_2D of inst : label is "6630C02930BE0AF816032C80000022201C4494D986E1423C01400661541851C6";
    attribute INIT_2E of inst : label is "D85B0BC026196C1996D96208B1D2E619471CCD8300DB7343D009C6E140666666";
    attribute INIT_2F of inst : label is "8252A00C2110318C2BFE46DA49B6926DA49B69273920010A13830ACD55000100";
    attribute INIT_30 of inst : label is "BE1D5F7FBE5D59757DB6F9757DB6F9756DB0F6DF0FB1F5BE5F63F49FCFFCFFCE";
    attribute INIT_31 of inst : label is "0483102C0968161208210A8001376472157CBCF9756532EAD801B0EEDB1D5F7F";
    attribute INIT_32 of inst : label is "7EB0A356ED02C33346C533346C132346C1007FFC80A8541C0830720581410008";
    attribute INIT_33 of inst : label is "8A161201E8A40E2DDAF2280B9F8BFDAA844AE7A80001032B93F208004AFAA121";
    attribute INIT_34 of inst : label is "2EA002002EA010412EA4921EC820023E8008007E93F9FF9FF9DE222C584AAF88";
    attribute INIT_35 of inst : label is "222A802A8022000000032417832EA4A25D4000001ECB23A8200003A800000BA9";
    attribute INIT_36 of inst : label is "FD5D75D75805D77775F777602AAAAAAAA00AAAAA8000000000000000000AAAAA";
    attribute INIT_37 of inst : label is "81E00A0000000101A54A0852A07367204028041A93FF014810000448240F775D";
    attribute INIT_38 of inst : label is "806018060180601810FF2036008A207FD0DC47FD00047FD00440611FF4289145";
    attribute INIT_39 of inst : label is "003C01200300702380040060300018000484062404044A080890100800030201";
    attribute INIT_3A of inst : label is "9E8E38E000000000000001044240000000000000000007C601C100FCE0360008";
    attribute INIT_3B of inst : label is "EB08CA855ABF414CC610E103A7B442A02D0800010949070DB041FF445295A4DC";
    attribute INIT_3C of inst : label is "4CD55FB37FFFFE0000002100AB105404A9068A59522211CFFFFFFC488AC2348C";
    attribute INIT_3D of inst : label is "980BC9B02F26C0B49341B1E30E6E0DE3C7873706F1C3C0608A214F06250A94B7";
    attribute INIT_3E of inst : label is "30E1330A5847BE200036C9B653810B9056FA66AE868200CC4444932850EBF294";
    attribute INIT_3F of inst : label is "CC179040A52242C43B888C18B10E622304492048B28921442D004C821894C008";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "B20134582600000000000000000004908652C0C0000000190072B694F0F86A85";
    attribute INIT_01 of inst : label is "6760EE079650964DC0DB292003390C0784C00800001320AD174524C14A42E4A2";
    attribute INIT_02 of inst : label is "3855372D9CC38C3050996B0D32C0D300D344258DCE6380700E1135A154C1E399";
    attribute INIT_03 of inst : label is "DB34D92669B24D50285842DE83331112CCD44416148281A2412126466A8D9057";
    attribute INIT_04 of inst : label is "5679783680B9A69B6DA469A6DB6936DA469B36DA4499A6C9334D36DB48D34DB6";
    attribute INIT_05 of inst : label is "A050405910C0B8021B9ADD60201A4403441114E69CD39904900800A44189CD8E";
    attribute INIT_06 of inst : label is "DB6CD36499A6C9355249E6489259998DAD94D3ACE45DB6E90992B822F0020038";
    attribute INIT_07 of inst : label is "2C60C0C20E19E0734D36DB48D34DB6D26DB489334D92669B24CD34DB6D234D36";
    attribute INIT_08 of inst : label is "0900010EC52220C988924822B29D225C12A8AA007CA80903098D8D8D8C022A16";
    attribute INIT_09 of inst : label is "1927113791141931648953092492491496745294C139965842400924B330A080";
    attribute INIT_0A of inst : label is "CB299ACB6618325AE4C8728019993221313CCCAD6D860C60C37042886DB28033";
    attribute INIT_0B of inst : label is "2D2B4AC8590C812904094ECB640948204A765B244A512253B2D9225289129D96";
    attribute INIT_0C of inst : label is "5B5B5927ACB698748C366D2B214B6B6924F196D30E8588ACEB58975AD4AB04B4";
    attribute INIT_0D of inst : label is "6D30E8D25B4C3A4B186CDA56425B5B59278CB698741A12DCC3E0B061B3611948";
    attribute INIT_0E of inst : label is "0484AB11A1D21B5B69C1836AAAC33259306C9364E30020644AC52AC9ADAC93D9";
    attribute INIT_0F of inst : label is "1128E180809889C1C0809A29A29A29A2B284D4D4D07B7F45B000000000000000";
    attribute INIT_10 of inst : label is "DBB3C96D30E9670A40B10B42C0B3B3B676CEDAC690A48009284AD2012C2A4893";
    attribute INIT_11 of inst : label is "C592DA615ACC141B76D6792D86DF2C96D30AD66080DBB3C96C36F167084C924C";
    attribute INIT_12 of inst : label is "D6B33262C99609A68C82A8022A960000000000006176D22C8B21B76D67B2D0DB";
    attribute INIT_13 of inst : label is "262644A93811E87468842E4188A002400A51A64D193808C242404042424240C0";
    attribute INIT_14 of inst : label is "D0A4A149429285250A4A1492009349285250A4A14942928525080449A5BB6CD9";
    attribute INIT_15 of inst : label is "B556AAC3A9322222448912232524964AB6C58333423211D946CAC2C4F50B9162";
    attribute INIT_16 of inst : label is "54D6D2952A54A552A9089C2274AC912D00934099332544A8C9992492291155AA";
    attribute INIT_17 of inst : label is "4160B650582D94160B610582D902C81CA5D8343836D936D936D836D8D54A54AA";
    attribute INIT_18 of inst : label is "0608806194200020F048482FC00B68082E1212D4AAAD264C8E4C891C995602D0";
    attribute INIT_19 of inst : label is "52936CD6CDBA016AADC94AB1C99EDC310162282D1C326C0B0520A51F50814829";
    attribute INIT_1A of inst : label is "6D436D437E86DAA64444444444DB6DB6DB48244326CB30D8204A5252B3516689";
    attribute INIT_1B of inst : label is "1B6216C290948CD9EDDACE1864D926190216C29094ACC8E4C2D2956956B48943";
    attribute INIT_1C of inst : label is "D9661B6216C290148CD9EDDACE1864D9661B4216C290148CD9EDDACE1864D966";
    attribute INIT_1D of inst : label is "945A241649271548B06F0B830B5C0C330C9B300A0000F5045510242D104E1864";
    attribute INIT_1E of inst : label is "D52A495AD3102D5C6DB25115C1071616D97B3496D916D92C9212492B78912238";
    attribute INIT_1F of inst : label is "8152332B014A76BC076C76C76CE59635F759CB2C6BEEB39658D7DD672C91AFBA";
    attribute INIT_20 of inst : label is "62B68C75959A960A00020C00428D101D9203484570090111546EA957556A21C3";
    attribute INIT_21 of inst : label is "B7296FA60DD86C96232ABCA6522530369ED3C2D94DD61EC32480486ECEF2A934";
    attribute INIT_22 of inst : label is "EC78849660A69F6E521BE9FC7CB27870BBDDE41427FDDF12405FF76C4BBD189B";
    attribute INIT_23 of inst : label is "610DE976B3721954D3104AA52424000000000000000000000000100CA4E52244";
    attribute INIT_24 of inst : label is "85188E02AB6888CE77A7AD9AD63449B22331CC05AD6B0137D26B8E0EC0C22C05";
    attribute INIT_25 of inst : label is "359E49B59ACF34DA49679A8E6398E534D366C0AC4DAC967922D8493109221849";
    attribute INIT_26 of inst : label is "42EB4BAC3711688352D99844650428924946592C2D824DAC967926D64B3C936B";
    attribute INIT_27 of inst : label is "54966F33994BB1BC5E56966F336D8DE2F2B4B319CD499C5E336A5C362DCCB6B7";
    attribute INIT_28 of inst : label is "74C44269B8C9BCCE966E326F33B59B8C9BCCED666326733A59BCD4C63131BC5E";
    attribute INIT_29 of inst : label is "581C29247039669918CEF19753464B4BF1ED62F5DD1A48C96E705B9ACDE7ED98";
    attribute INIT_2A of inst : label is "C0CC0070C5C152201B608C30229411B6FECDBD95270E46311903BB0A121440C1";
    attribute INIT_2B of inst : label is "970725D5ABEAA72DC0EE1076BDF0AE1D410426F530AB853210314000000A4C76";
    attribute INIT_2C of inst : label is "8CB8D28654D9432A6C24F42457F614FC3CD89049D5207A2C4A056E6A815736B9";
    attribute INIT_2D of inst : label is "44AEB60AA527569D142A0958000057D7FC2D288134A706AC57CEA338DB8E36E3";
    attribute INIT_2E of inst : label is "985B0BA074D04951049041802530B592D4D2892A40925AE0240974A702666644";
    attribute INIT_2F of inst : label is "0259DB2CB311AD6347FE44969125A44969125A45AA40024C9292488AAAAAABFE";
    attribute INIT_30 of inst : label is "BED19F7FBE919A467DB6FA467DB6FA446DB694DF6FB539BE9F6F392C00000000";
    attribute INIT_31 of inst : label is "CE97116CD84D35B2C218CC8801232460067CBEFA4665B488D9FDB68CDB511F7F";
    attribute INIT_32 of inst : label is "7EFD3224EBC2D39356E338356E339356E3007FFC91964EBC0CB2E22D935B0020";
    attribute INIT_33 of inst : label is "35F9EFFFE28B31D66520A3F4607408220B2518500000CC946828807FA5052121";
    attribute INIT_34 of inst : label is "48CFB4DF48CBA69C488924D2938D74A637D3EDE725800000001EA0D367BD57A8";
    attribute INIT_35 of inst : label is "282AAA8000282AA002814B97DC48C8B4911B3FB6D2934A238FF5DA33EE77D232";
    attribute INIT_36 of inst : label is "F5D7D5FD5805FD7D7DD7D7C02A0A002AAAA00282AAA00282A82800AAAAA00280";
    attribute INIT_37 of inst : label is "ABEFF2A000000012010AA000AA000054054001400000A000A085400A8007D7F5";
    attribute INIT_38 of inst : label is "505415054150541505FE01700100048FC30148FC30548FC300480523F0C05201";
    attribute INIT_39 of inst : label is "45815608B02AF1400A005002802800140000280404500808A010114001400141";
    attribute INIT_3A of inst : label is "263618600000000000000100000200000000000000002F800BC005F0017000B0";
    attribute INIT_3B of inst : label is "494CE11E933FC970F820E2C9716E59A2DF000101070707079203FF446318C0BA";
    attribute INIT_3C of inst : label is "D0367EF4FFFFFEC6010842189B19B6658942B656E31DAD3FFFFFFD6112D765A6";
    attribute INIT_3D of inst : label is "1C1B81E06F07C1B09341B4EB5E6C0DC9972F3706F4CBD000150563842B0BB2DD";
    attribute INIT_3E of inst : label is "32E36CA6BCB13AB1003659B2CC42C5129B51B800000200CC555593695AE7E9B4";
    attribute INIT_3F of inst : label is "CD2308EDC0BB66E313883CD9B8C46207306DB26EE0ED98764D0082C010965938";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "0C324C0D6400000000000000000032C78612042000000004390BF10381213967";
    attribute INIT_01 of inst : label is "20682C004F80E13FB7208CB24884B4688D1C1800001CB23A3100D3AC11662098";
    attribute INIT_02 of inst : label is "DCC66D9B75AEA1B706F6D6B9658B965B963287498118809482026EDE518142C8";
    attribute INIT_03 of inst : label is "DB34D92669B24D5AD4CC66133999CCCC6663332C5ECBDE1B6D8D9BB3243A6846";
    attribute INIT_04 of inst : label is "0D0EC65B4039A69B6DA669A6DB6936DA669B36DA6499A6C9334D36DB4CD34DB6";
    attribute INIT_05 of inst : label is "10C2DA0C26189481656322926CB50D969256E308610C25B2CB24920B26E06361";
    attribute INIT_06 of inst : label is "DB6CD36499A6C935692431A1993438AB12F28C1389330D9E6CCCE60388E2803A";
    attribute INIT_07 of inst : label is "1F56834EA8634FF34D36DB4CD34DB6D26DB4C9334D92669B24CD34DB6D334D36";
    attribute INIT_08 of inst : label is "64B64C66A48F872719924838094449338828AAAB2A000025128707070462AD9B";
    attribute INIT_09 of inst : label is "0E9183C843C0E4E310491849249249C34D1B08C313244181A6596096088602CB";
    attribute INIT_0A of inst : label is "2084E1B082C8D9A656DB9919C5C68986CEC216C80A61981980CCB863DA40498E";
    attribute INIT_0B of inst : label is "51B46D246C24588462C421B082442112210D84162118B1086C20910844884361";
    attribute INIT_0C of inst : label is "642424103E484322E19990A78D6C84848203C908644A6253A02769010610F746";
    attribute INIT_0D of inst : label is "9086470B2421916CC333235F1B642424101E4843226059221956C30CCC8D7C29";
    attribute INIT_0E of inst : label is "137B12C30D2824904D2EC8C223BC29248912CC831E6D93997539C4361212083C";
    attribute INIT_0F of inst : label is "ACD8E2C2CB666E1C6C82E3CF38E3CF38620707070C84E4CC7000000000000000";
    attribute INIT_10 of inst : label is "24482C9086469C2154C14C0314CC4C418831053146534B2493250925D0CD0F0C";
    attribute INIT_11 of inst : label is "1A59210CA5384664890905921521D2C9086529D23324482C90A90E9D23B24933";
    attribute INIT_12 of inst : label is "094ECD302740C61CB328000280180001FFFFFFFEBE892C6301C64890907922A4";
    attribute INIT_13 of inst : label is "1D71303498664BCDE4449A8DF7D50B8C2D22D138669351189898989A9A9A9A1A";
    attribute INIT_14 of inst : label is "1B33346468C8D191A3234649034E6CCD991A32346468C8D191A013A75A6699A4";
    attribute INIT_15 of inst : label is "CBB9770A45A189891224488580B20030E1302E11210C4C4C5A631A30100C828D";
    attribute INIT_16 of inst : label is "1644C0DE0B231188C49006401DE348B180CB63588CD23446C46696DB059EEE5D";
    attribute INIT_17 of inst : label is "8C060863018218C060863018248513E2DA28C848E821E821E821E82471037831";
    attribute INIT_18 of inst : label is "2857909247BDEF8F496163909EE401E1C258590208329D2377B336EF662C1B98";
    attribute INIT_19 of inst : label is "294E1B80B36166C0DA6CA4266440A18225644CADA19991A4758EB0A7665D63AC";
    attribute INIT_1A of inst : label is "8064806484C90178222222233B2492492433B09999248664202B095859ED9C14";
    attribute INIT_1B of inst : label is "CCB2110AC2D636377B3530C3332490CC92110AC2D636377B1D294294294A1464";
    attribute INIT_1C of inst : label is "2490CC92110AC2D636377B3530C3332490CC92110AC2D636377B3530C3332490";
    attribute INIT_1D of inst : label is "C00018450491C0912349F47CF7ABF3CCFF66CFFFFFFFF7FFEAC0909847F0C333";
    attribute INIT_1E of inst : label is "298B0C6B1B42E830082B7C49340AC0C4903A82400645140061C124129144880D";
    attribute INIT_1F of inst : label is "C1CC45060EB1A849BC18C18C1B32C9C628A665938C514CCB2718A299964E3145";
    attribute INIT_20 of inst : label is "9548529A4A61492A99B9B8ADCB07A6AA2E6A37206E0FB0AAAA5DFAAEABACE5CB";
    attribute INIT_21 of inst : label is "739490581CC9DB600114147B2872C249612C27243219612C9249A19030514CC2";
    attribute INIT_22 of inst : label is "2187334991B840E72864162A06490CD9CCCC903984CCCDC9249333272993CB60";
    attribute INIT_23 of inst : label is "CC10F4643A351ACB1896C0C200C0000000000000000000000002000C80A4050E";
    attribute INIT_24 of inst : label is "41DF448C03F6E37398C918AE731D2DDE298C340A52944CC804B235447798191A";
    attribute INIT_25 of inst : label is "9241264249209321209041694AD696C96C9744523212090459896DC92DBD096E";
    attribute INIT_26 of inst : label is "43824E396CDCB6866BA6712310B2964934390412125C32120904590904820C84";
    attribute INIT_27 of inst : label is "092D91C99924464720096D91C916323900596CE472E6472000C358E4DA28E4E8";
    attribute INIT_28 of inst : label is "298361C6432647206990C991C80A6432647206990C991C81A6472E1C9C464720";
    attribute INIT_29 of inst : label is "72766EB6A9421966F7B7DEEF8F78B434AED19F0D62E3679692A962633239F6C7";
    attribute INIT_2A of inst : label is "A03A090C2040719830C218110E08404983832938B09135AD76DDB0F4844E9393";
    attribute INIT_2B of inst : label is "4886871CE35578BA20798C3DE491FA17AC13B21D06089289CFB400000065200D";
    attribute INIT_2C of inst : label is "E6466D73AA46B9D524523CBC9CBA26302C799B3624503CB6405062B81471C845";
    attribute INIT_2D of inst : label is "2330DB20B1B846E1160B6C60000002B68C15B64987910B3F2165788E65639958";
    attribute INIT_2E of inst : label is "D85B0B9036596C5D96D9665DBD96F6D9421C458B42DB7BA0748987910C222222";
    attribute INIT_2F of inst : label is "392D1616D8EEE731D3FF76DADDB6B76DADDB6B773B7FFE64CB5B60ED55555402";
    attribute INIT_30 of inst : label is "BEDDDF7FBEDDDB777DB6FB777DB6FB776DB6F6DF6FB5FDBEDF6FFDBFFFFFFFFE";
    attribute INIT_31 of inst : label is "78ECEED63321E06B6CF073240C8DD121177DBEFB776DB6EEDBFDB6EEDB5DDF7F";
    attribute INIT_32 of inst : label is "0190CDBB393C2C5C2819C5C2819C4C2819007FFEDEEB2966125D8DDADE060093";
    attribute INIT_33 of inst : label is "8007FDFFE8A0C7799F8228019FDFE088B09AE7A80000306B862888001AFAA121";
    attribute INIT_34 of inst : label is "6EEFB6DF6EEFB6DF6EEDB6DEDBEDF6BFB7DBEDFFB7FFFFFFFFDE82009FF7FFA0";
    attribute INIT_35 of inst : label is "7FD55555557FD55557FB6FB7DF6EEDB6DDDB7FB6DEDB6BBBEFF7DBBBEFF7DBBB";
    attribute INIT_36 of inst : label is "002880AAA008AA802A02A8007FF5557FFFFFFD57FFFFFD57FFD555FFD55557FD";
    attribute INIT_37 of inst : label is "0010081FFFFFFC01FEF01FFF01FFFF43F03FF03FF0001FF81C703FE07FE802AA";
    attribute INIT_38 of inst : label is "00000010240902400001F40FF8FFF07010FE47010FA47010FF47F91C043F91FE";
    attribute INIT_39 of inst : label is "907E41F20FC8003F81FC0FE07E07FF03FFFE07FBF80FF7F01FEFE03FF03FF000";
    attribute INIT_3A of inst : label is "4140C308000000000000010000020000000000000000007FA03FD00FF40FFA0F";
    attribute INIT_3B of inst : label is "B433234FFC9F1480FE40F8844A496D101501000205010D059501FF3318C6378E";
    attribute INIT_3C of inst : label is "407F4891FFFFFF6300C6118CD0E42912ECBC05808CD1192FFFFFFDA24D0CDA19";
    attribute INIT_3D of inst : label is "F20C2F0831BC60CEDE20CA36A1C106146C50E1831A36663DBA9CB001929659F5";
    attribute INIT_3E of inst : label is "DD9B7A86B862F70C00ED3769BCC1A6EC3257A8000001015044477E84B0D3ED42";
    attribute INIT_3F of inst : label is "84CB07831FEEDC3ECE7662370FA39D9883DB61DB9DBB70CD1801372CA6C9340C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "1413047612000000000000000000328786024220000000042521692B218B73B3";
    attribute INIT_01 of inst : label is "226868002E80823F9A900D92D91FBC018405440000081E2A2000E02807641010";
    attribute INIT_02 of inst : label is "5FA680C0402805A6068310A1041A105A10620C6A75918C3116208207053E1C28";
    attribute INIT_03 of inst : label is "92A695B54D2B695AA0C46275B111888C44622370CA594AD925050AA002212004";
    attribute INIT_04 of inst : label is "002F4EC94D2534D249354D34924DA49354D2A49356D534ADAA69A4926A9A6924";
    attribute INIT_05 of inst : label is "3C713032458800804502175624440488D2DA220440881492DB2496122E402540";
    attribute INIT_06 of inst : label is "924A9A56D534ADA5600097809000A47813D385361B0410362440820218154958";
    attribute INIT_07 of inst : label is "40F5018C50A4E44A69A4926A9A69249B4926ADAA695B54D2B6A9A69249AA69A4";
    attribute INIT_08 of inst : label is "64964C67A40D0D4008924830010C000390A82222800000070B8D8D8D8C010345";
    attribute INIT_09 of inst : label is "0E0081A50181A80100C9104924924981001E0087312C820FA2484094100C024B";
    attribute INIT_0A of inst : label is "818CD0D142D851D65249111B850601025A5017783AD348348104F1454920695B";
    attribute INIT_0B of inst : label is "68BA2E846824588C62C460D142C4631623068A1223089118345091184488C1A2";
    attribute INIT_0C of inst : label is "5200000034000222C11100E50D6A400000068000445D516A01052008041873A2";
    attribute INIT_0D of inst : label is "0004468E0001116A822201CA1B5200000034000222D0F0041152A6088807282B";
    attribute INIT_0E of inst : label is "1B691E8B1F7422F1CF66D94222B464925B2A8A411B25508B56A9461500000028";
    attribute INIT_0F of inst : label is "E488E2C66A07E5186482410414410414600282828C44A4DCB000000000000000";
    attribute INIT_10 of inst : label is "928038000456560554A40A0294AA2A21442886A382605F6593269B6CE9EC2D05";
    attribute INIT_11 of inst : label is "9970000894AE0A52500007001C95CB800044A5705292803800E4AE5605EADB6A";
    attribute INIT_12 of inst : label is "852B44084015C51611000002AA940000000000009A54A4250145250000500392";
    attribute INIT_13 of inst : label is "16A8A838551A0672BBAA6924C0E00120362E402D221310989898989A9A9A9A9A";
    attribute INIT_14 of inst : label is "8D191830306060C0C1818301018066468C0C181830306060C0C002C05D6F5BD2";
    attribute INIT_15 of inst : label is "8110220EFCE111102040810601A00210A2A0FE00001478844C220C4025588346";
    attribute INIT_16 of inst : label is "1444C0CE0A231188C4B88AE229450890C08A31508862344684431249048C4408";
    attribute INIT_17 of inst : label is "D82C14360B050D82C14360B0508693D049702C23B050B050B050B052B1033831";
    attribute INIT_18 of inst : label is "2047D01006B5AD0C794141028A40034304505086410100804200108400340A8B";
    attribute INIT_19 of inst : label is "A18A2A83A12FBF44687E8064448381066D4CC5A8811100803506A087E44D41A8";
    attribute INIT_1A of inst : label is "0060006014C001F422222222295249249213A99110000444206A195061C6D450";
    attribute INIT_1B of inst : label is "8892128A82D438042006A08222000088D2129A86541804200EA1035035A91860";
    attribute INIT_1C of inst : label is "000088B2128A82D438042006A08222000088B2129A865418042006A082220000";
    attribute INIT_1D of inst : label is "840A08083001A1F3E7DBFFABFCD4FD7760BD1AF55C30FBC44000008D03E08222";
    attribute INIT_1E of inst : label is "ADC38C6B1A01D81E38E1388F580C828DB036510452087045228C001653881010";
    attribute INIT_1F of inst : label is "8084540A08000001B52852852A02810425D40502084BA80A041097501408212E";
    attribute INIT_20 of inst : label is "49A4691D0D518540F606F1C21C022C77181193604607802AAA1172A8AAC4CC99";
    attribute INIT_21 of inst : label is "51104850088949211000146A20228249412822006949412892498148210008A3";
    attribute INIT_22 of inst : label is "6905210910B400E62052142A2C402C588888821B10888C8924C2222221128804";
    attribute INIT_23 of inst : label is "C800D06423341ECA4C82A0F398D8000000000000000000000002003C01200C04";
    attribute INIT_24 of inst : label is "40D504C00263D3D6B18118B8D6B42D76098E380C631868EA0D9E71603F903980";
    attribute INIT_25 of inst : label is "1000240008000200000001294AD6B6496D95C01220000000D089248924910925";
    attribute INIT_26 of inst : label is "400240A120D296802A06D8062092440010F00042001420000000D00000004800";
    attribute INIT_27 of inst : label is "113500816600C4020013750081022010008BA840204402000147088402080408";
    attribute INIT_28 of inst : label is "2B0125440204020075008100801D40204020035008100800D402041618440200";
    attribute INIT_29 of inst : label is "33272692A887094216C7D88FAE20B810A8C1020902C1279302A882422011F2C6";
    attribute INIT_2A of inst : label is "906908A420807198114008308E0C20CC02204238A08114A55A14201484029919";
    attribute INIT_2B of inst : label is "0086071C630030A020608431C001F0032003A20D0F090001AE80000000568450";
    attribute INIT_2C of inst : label is "D545342AA90A155564422C9C89DA22220C399A22AC6030A6401061B804708005";
    attribute INIT_2D of inst : label is "23925B60909A446902092448000028160C3096489392839EA014354D56535514";
    attribute INIT_2E of inst : label is "48090180120B2448B24B3659948652CB02484489404929E07400939286222222";
    attribute INIT_2F of inst : label is "7027721648678D6B43FF32484C92132484C92132113FFE54A959506400000002";
    attribute INIT_30 of inst : label is "BEDDDF7FBEDDDB777DB6FB777DB6FB776DB6F2DF6FB5FDBEDF6FFDBFFFFFFFFE";
    attribute INIT_31 of inst : label is "6A74EF525295A0A974D8637408144205177DBEFB776DB6EEDBFDB6EAC35DDF7F";
    attribute INIT_32 of inst : label is "01A045A139342ACA3431ACA3431ACA3431007FFE4AA93BA616DE8CEA5A0A00F3";
    attribute INIT_33 of inst : label is "8A1A1201EA8C0CAEEAAAA20A212A002804600800000103803800000060002121";
    attribute INIT_34 of inst : label is "6EEFB6DF6EEFB6DF6EEDB6DC5BEDF6BFB7DBEDFFB7FFFFFFFFDEA22C684AAFA8";
    attribute INIT_35 of inst : label is "2AAAAAAAAA802AAAA8036FB7DF6EEDB6DDDB7FB6DC586BBBEFF7DBBBEFF7DBBB";
    attribute INIT_36 of inst : label is "AA8000AAA81200002AA800000000002AA000000280000002800000AAAAAAA800";
    attribute INIT_37 of inst : label is "340003400000014400034000340000680A8006800400400343028015001802AA";
    attribute INIT_38 of inst : label is "AF2BCAE298A6298ACA000680060007000C003000C043000C003000C003000C00";
    attribute INIT_39 of inst : label is "0A002801400502801400A005005000280000500000A0000140000280028002BC";
    attribute INIT_3A of inst : label is "60204000000000000000000000000000000000000000500034001A0006800340";
    attribute INIT_3B of inst : label is "8215602FF51FD9FF0080F180DEDB37107404000804000C048C00FFFF0842178D";
    attribute INIT_3C of inst : label is "007F0001FFFFFF610046118CF06CEB22E8B41C838DF30D6FFFFFFDE00085410A";
    attribute INIT_3D of inst : label is "D6087D5820F5208FEA208C3AD343043874E9A0820C3A3A04B054E0011ED261E0";
    attribute INIT_3E of inst : label is "CE9A6E15B030D78800849424BCC0C66032578802AAAD011444455A469083E723";
    attribute INIT_3F of inst : label is "94DA06A53EAA541B0472225506C18C809F49214A8CA9584508012224268B1006";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
