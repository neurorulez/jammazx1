-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity bangpcm is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of bangpcm is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "57683C05B777A04A4DF9278D76EF901E848DE740A847BEDF3100B05C8329F7FE";
    attribute INIT_01 of inst : label is "F4ABF734608CC6AF81EA08335F080578BDCDA5E1F9E459D32AED893BF046E148";
    attribute INIT_02 of inst : label is "89E08A07F3341AA6DDE3F3579665B6B521B8B31BF7BF49582C090423727DBA47";
    attribute INIT_03 of inst : label is "FD8E5176EB3D2552AA4B344082FE5CB9940AEDCA1D836BAD3BCC382FCBABA25D";
    attribute INIT_04 of inst : label is "1AAF67A8D61FA6CB9484827D36F0A40551EAC04B8D5B3EC59A2D306D29917750";
    attribute INIT_05 of inst : label is "1D9FE79254C1862DB6783D7AA4DB76CD2EB1B96A3443C7A37AD966A28B1F2A19";
    attribute INIT_06 of inst : label is "D96F64E1B1C7821BA6612A87FDD185181CAB6D7A6472201DB128BFC1C72C6250";
    attribute INIT_07 of inst : label is "1EEAB44E1880690D46BB6E4B1052585E9E4667DC4D890D7A186CAE82586B5345";
    attribute INIT_08 of inst : label is "D93D797271E880A372681E768ED8BE82ABC6E21A6745CA184813DAF2CA151FF2";
    attribute INIT_09 of inst : label is "411E46C58288BFE8A722EE9DB0F1034DF90CB3A498A7D28F123FF2BAA7B7897F";
    attribute INIT_0A of inst : label is "C848145D3EAA56F9D177D525C770D036096F27E0B9B0812C3805FDEA8FE96F29";
    attribute INIT_0B of inst : label is "C769D284DB1F04D63E37D564567F5B47BE72D6F8122E16C726FF071DF6157684";
    attribute INIT_0C of inst : label is "A7434C32668B215FCFE478D66EFA45A7559CDBCA226AEE368548E4F9E5479684";
    attribute INIT_0D of inst : label is "EC03ED1CD03B657F933546B989387DBCE5F4C0FC9FF0B2E151C54C74C6209D29";
    attribute INIT_0E of inst : label is "69063DA2DAB43EBE685A30F6F55550CDDF31083B2119DDDA9E95A5B41190A5D8";
    attribute INIT_0F of inst : label is "2E20E2752538D86425BC04506FCD6466BF9DEE81BBAEF580D3FD5F4F8A39D6A2";
    attribute INIT_10 of inst : label is "8F836307E8AA90282023B933EF38C35EF186FED775C0CD14A83BDF4764CA5120";
    attribute INIT_11 of inst : label is "DBB8B76E51716E67668B6FA0D7B8F831276242BB9B5FADC851C28E904BCC7E3B";
    attribute INIT_12 of inst : label is "33DA63D3FF83DED313281E1606C9DFDAEA660C806DC2431A8750E4DED0B6EFA9";
    attribute INIT_13 of inst : label is "04364466E574AAC0697D395FF38C2D31510E1442049828F4121B31FD01DA7F6C";
    attribute INIT_14 of inst : label is "9DFF5094CF1C131753D0D6FCECB78FE92E349232EE74A7F741CBBAB230A2A4CB";
    attribute INIT_15 of inst : label is "B2AC7E33E228513A2D4DBFCF17309FADE55FECB4E265986CEA36F98C2F658ED8";
    attribute INIT_16 of inst : label is "37EEF978CCEE284E4358C77591F319AEF3A210337B7A2F40141593AC55B3FB02";
    attribute INIT_17 of inst : label is "B1CB72108147E74136BDA4A6915160B8A3376991A866CA1A57DD93699242DA9E";
    attribute INIT_18 of inst : label is "173002D64BA213AAFE8DD48660348ED39E6B2FE2A67550A9569A24451B878A6C";
    attribute INIT_19 of inst : label is "FFC64872A3CC6AF31B8CB7DBCA4561C169978EC7CE02C04046C92E9C98629A2A";
    attribute INIT_1A of inst : label is "35E85E011C25F796E2333F95E3FA468B1BAADE69EC172D8B1F69D35268326113";
    attribute INIT_1B of inst : label is "2FC8197B708B6ECB6E5A0B0EB8D52747ACEEB1BCA9F084874EE670A3B9A282F0";
    attribute INIT_1C of inst : label is "E8C463C14320AE5319D870D6B2EC9C2AF51EFD928400AD8E0D93F489BD845968";
    attribute INIT_1D of inst : label is "880F145D4A4A374B883405A68AAF555EBEBBB22CA43EE1D42B4420B4A25939C6";
    attribute INIT_1E of inst : label is "34A80E093F286ABEA878AD6AC40843514CC94C8EF43CBF2C4430EE2972B4C4A7";
    attribute INIT_1F of inst : label is "015B795556B4330FBD5E1A00A3A7364EFBCD430CD4CD21C81453119C3CA4A72F";
    attribute INIT_20 of inst : label is "833D1E1CBD58D17BC9FE68F681AEBBBC81CC4A415BBAD854A5C3A70545730800";
    attribute INIT_21 of inst : label is "297C709DA5ACEF2DDCF4B7D09B894E56AE5472C813BFEE10DE299F357F23FDAA";
    attribute INIT_22 of inst : label is "60501990DD1C0FC081E74E31E42F4AF72B158D51373B52F993A5948FC17AFF35";
    attribute INIT_23 of inst : label is "3302E0166E6139F11CA99E5CB4E6003380E4F502BC126BC6BCC5BEF3D16A174D";
    attribute INIT_24 of inst : label is "84607E17C43639FA03984FF78C38CD8206072E7D4431E779FB9D48D15EA2C387";
    attribute INIT_25 of inst : label is "0FF3E0001FF10400060FFFF81C73773181C41980E46E0CDE7E0C6079CE640101";
    attribute INIT_26 of inst : label is "01F031CE78C6E18FE0CFF1C70078030730664A79A5200E663EF8C7FE31831F0C";
    attribute INIT_27 of inst : label is "FFE3DE07C7FFFFFFF1C183FF1EFC3C3E4F8701F80FFF80FE00F8063E0701FF80";
    attribute INIT_28 of inst : label is "DF00001FFFE007F807F801FE00FF801FF00FF001FFFFFC000607FFFFFFC0000F";
    attribute INIT_29 of inst : label is "000000003FFFF00000001FFFF0000F180003FFF800FFC1E003E703FFC780073F";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "24A4BD82D0B8186E78D3E2A9823EB642C5C0ADAA61FB1764F7CA706F4A4E1E56";
    attribute INIT_01 of inst : label is "657E35F52911DEBB719F72D376961D57EE13911BCD133860FFAE763B6A69F831";
    attribute INIT_02 of inst : label is "0FE6066CCFF7041509E97103051DEEB88F9BBDAE11E7A1DBE169F97CE47D29A2";
    attribute INIT_03 of inst : label is "8656C7996EFCE3231F9F3C69E990AD8C78C67149CE70F4DA6CDB153039C9A609";
    attribute INIT_04 of inst : label is "2B03BB97369E57731D07FAAF22C0DA4EC7F3A9B59F307A050809C66D2BD99B62";
    attribute INIT_05 of inst : label is "F5E2DD13F3EA005758062E1D328B53FA22ADA7BB3A3C046C3B3823DA957E1A8C";
    attribute INIT_06 of inst : label is "91CED50C38C040F9C465BCE53855C4D98CC8768341F1B1A274E6F0061EFF9B82";
    attribute INIT_07 of inst : label is "104EB4BD5983C1650B510A58F2C5FBC7857238D214176A48CAF779D8966B0AE3";
    attribute INIT_08 of inst : label is "5D8DBC5372ABE5642029A22C86ACEC90060577B771283869535B145742D01500";
    attribute INIT_09 of inst : label is "CC30BEE7087CEF8D0402AC2D047561D93DA85D3EEB9E538F2F3B6057DE9193D2";
    attribute INIT_0A of inst : label is "24683B312611B9D7F6E1965CCA2105A8B9F22FBE5858EEEDDD290BA817D7D604";
    attribute INIT_0B of inst : label is "E6063226EE346309559480976711726047D5F5905AFF6B4F6A4174AC6D5A02AA";
    attribute INIT_0C of inst : label is "5AE0BC4C37E92F8969D421B4D5F5942AA69C93F3333FFE4E6C91AFA22AA45E60";
    attribute INIT_0D of inst : label is "9B55BCB3CC2D2EE34E087436C6FC46293C3E5D6FCD5511D4843709ECCB664B4E";
    attribute INIT_0E of inst : label is "07FDB45A9A5A3A7EAF895A08093C2C75D8786BCACBC49731A704605540F7D342";
    attribute INIT_0F of inst : label is "5A9954200C01CD62A7C81B64E62A677784EAFF646D806012282C610147D46ACB";
    attribute INIT_10 of inst : label is "2EEF60D6670AB9BA4A765FFC4C1E49D5DDE63D6F5C6EFEE744ADB38B15BE07BA";
    attribute INIT_11 of inst : label is "93ED162A9FEE018FFE4A14B2CEB789A6788761DC774AEF175D4530197481AA55";
    attribute INIT_12 of inst : label is "3B8D6BECF1BB608DE47AB9B3DB03210F8574D141DFA9D278FE2576BE6CB418D0";
    attribute INIT_13 of inst : label is "4210F5899D5D9ED102289A402169269502F323AAD688990F792CE7997A44ADD2";
    attribute INIT_14 of inst : label is "EAC7EBFB810E3F187F21EA44C77021CF3B526C2CA1EC4FF25C9158E1CFC2CD47";
    attribute INIT_15 of inst : label is "62F6BB76B54966B28673AD3A2977B4D8E826A1AEF76CCFA5C8B1EE842C493FBA";
    attribute INIT_16 of inst : label is "E6FB82B9904BACE40416F2FBA8F9BB64F6653D12DE410B4AB0480B1AEC6A19DD";
    attribute INIT_17 of inst : label is "C057B3172524EBA566D0177DAE21E96ABF043D2B2F0FAE3F65630FEA5E39EDC4";
    attribute INIT_18 of inst : label is "271A8F3491E06DEEB422A3C3249F8717E8CE021650DC8A38F1891328B5025942";
    attribute INIT_19 of inst : label is "91F76D1AB6A57B31B29EFD8FD3A7574BA273C853E6018659160A4E3D89713A13";
    attribute INIT_1A of inst : label is "61744E8E4F32210B10AF2E81EBD525F569871AD8185061638E2DEDD9C02FC0AE";
    attribute INIT_1B of inst : label is "503AA5658976EC057E2C09D7BD8F3FD2CDCA91DBC32CB1240804753EC75854DC";
    attribute INIT_1C of inst : label is "DCA0B426D59E1B5CF14B18FD2A4FB94E42E90FE1365E4604282F1EE971B25BA1";
    attribute INIT_1D of inst : label is "A1960DBCDFD50EF92AF9B0D073F538DE6B563A5C63FF5385826F4E16A66AB9A9";
    attribute INIT_1E of inst : label is "C5437E0E3FF41AD7ABFB8F2CE1F4C220AB569357D8E2956393B2DE3455989291";
    attribute INIT_1F of inst : label is "01990193DB721CFF8B3BF92F92FEDDA8A6ECD29002EB34E43933D7DD7F35B832";
    attribute INIT_20 of inst : label is "08C311FC11199B02F1FB98F58435C08381F87B4534321A5CCE386F0B9C54D800";
    attribute INIT_21 of inst : label is "0F1E710379881B339EF3101FBC7971CF35CF81FAAD6AB15A404E1F3900E001CE";
    attribute INIT_22 of inst : label is "E06007E71CFC0FFCF1E0CE21CBA719FA330C8E6E0CFC6101B043F10FC279FFE9";
    attribute INIT_23 of inst : label is "C0FE1FE67180F800FC31E06393F9FFC3FFFB0CFCC3F013C13C393EF6B1B3A724";
    attribute INIT_24 of inst : label is "FC000007F80E0603FF878FF863C00E01FE071FFE7BF1F81803E3271A6191C3E7";
    attribute INIT_25 of inst : label is "0003FFFFFFF10000060FFFF81C03F03F81FC0180047E00FFFE0FE0780E1801FF";
    attribute INIT_26 of inst : label is "01FFF0307F3E1E0FFFC001C7FFFFFF00F07873879CE00F87C007C0003E7F0000";
    attribute INIT_27 of inst : label is "FFE3DE0007FFFFFFF00183FFFEFC00000FF8FFF8000000FFFFF807FE0001FF80";
    attribute INIT_28 of inst : label is "DF00001FFFE007F807F801FE00FF801FF00FF001FFFFFC000607FFFFFFC0000F";
    attribute INIT_29 of inst : label is "000000003FFFF00000001FFFF0000F180003FFF800FFC1E003E703FFC780073F";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "0EB6B81A8D7C4122961AAF8B3FE0154EDA382F3348FD9FE73BD35AD949255B46";
    attribute INIT_01 of inst : label is "507A5F5F8DA803D4536A071464E305E55155274A681052B13D36046E73409BA7";
    attribute INIT_02 of inst : label is "46B4CB16964E745BA4844D694915B4151D296AF4DACDADD2B74FAB0B12D7A2F8";
    attribute INIT_03 of inst : label is "2B70A229C5204A533FE35424B02ECCD7ADEB4CCAB0DA83ECFD74641552C274A1";
    attribute INIT_04 of inst : label is "0EAA7FCA961541E0FA4E9575A078A3EC87D462DAE7E7A48AAA5B54D0EEF56D00";
    attribute INIT_05 of inst : label is "C9C659FF5406ABB2C957CA532EE56C90B91A9961A6AA7549BEAD7A742E129012";
    attribute INIT_06 of inst : label is "86A09BFCE56C8552D7CA25992C01B222BEE4076914A50A75342BEFD6C8519C99";
    attribute INIT_07 of inst : label is "5C964FE493ACD33B45478542A7922267DE31A632DEE9696F3EB08B17BF506274";
    attribute INIT_08 of inst : label is "08EBFA77B687AC739CE382611C390F80A3D045538E49928921F0A1640B2FE181";
    attribute INIT_09 of inst : label is "69B52BA9BB569C24C6E81A783CA7B79AA874C520DAD49B412F166BCF6656D0A1";
    attribute INIT_0A of inst : label is "B660803B30C19D09DB0A4CE948E8CFDCA797021FAC7004A4F4D379360D52A631";
    attribute INIT_0B of inst : label is "F8D2C23A4C62F4299C2152F46B1BDDB92D381EADF9991A3CB233FA56B77F528F";
    attribute INIT_0C of inst : label is "A239A8424B9681DEC4BE4F6A8B75951CC102F6891F555436A5B0D5AA033E7CB0";
    attribute INIT_0D of inst : label is "3D308F18A260A6D1F4D2ACAE15A5F165655D8892735A2747C34FF89151E94882";
    attribute INIT_0E of inst : label is "6CE6A1703E790B8F9052485109FB82592F671F7405C9F5C066A039C44A4D5DC9";
    attribute INIT_0F of inst : label is "D3D10D4D37DA8D5240991EF68B3E5A758248A056EB338EA7886E80CB1B4AB571";
    attribute INIT_10 of inst : label is "CE173013E062301C4FCEA52EF9DD91FA89B19E772F0013A5F2E0DEAD01C85942";
    attribute INIT_11 of inst : label is "0EE27BF688AC2747F7536B49992687BFE1AB9A5B816E0889F66154851DABE52F";
    attribute INIT_12 of inst : label is "2FF0CC0B71932AEB6E067C598E309E48155EF1961E8392F534171F9E293A506B";
    attribute INIT_13 of inst : label is "E40F42305196DF0FA2BCD108610E662C752C07B8226BD4AAE8815719F8D49D17";
    attribute INIT_14 of inst : label is "0DE4D0F4216A42C422B6A3ECEF4C0E229F8E0820CAB059446B3925E4B8BEAAFA";
    attribute INIT_15 of inst : label is "BF74C63CB59E7846EA3E6B394535AE05216E9EE6D7353AA089EE36951ADBB693";
    attribute INIT_16 of inst : label is "283EF5DFA689235BD64FDDFD50CD9DB7165481619F09DEA670B970A0B0D1988C";
    attribute INIT_17 of inst : label is "003300A035C8A0FC7703B2BD750579A8EA538499A5873F283E7F537F8177F20B";
    attribute INIT_18 of inst : label is "C91BDC0C75C94D394E027A7E8C0B4F84DE8EBC9C7A42542EC078F3CF9E48E1EF";
    attribute INIT_19 of inst : label is "7C73DB180CC9864652EAF0CB5B660D67A5F0C74FF4AAFDA305438E6E336BD043";
    attribute INIT_1A of inst : label is "CE6ED1A06D394E4408D740C9E6EBAB4E4384026D50391E4505BC9E76282DFB41";
    attribute INIT_1B of inst : label is "5FF99072062E1048AE1AB367AC0B4F8B0C4CB1E5F137A3CAF17E51C1AA1698CB";
    attribute INIT_1C of inst : label is "BF88983DCC80F81FF668770BCDDB3C71D5F2015F70C0A802343119B9A984B29E";
    attribute INIT_1D of inst : label is "609BFC23C3CE0087367E781BFC530161E6E42DC3E000600DA2F58E2D718D391A";
    attribute INIT_1E of inst : label is "FB0781F03FF806F06C0730EF03FDC3BFC84FBEE09F418CE01ACE41C39874E48E";
    attribute INIT_1F of inst : label is "01E701EF23F1DFFF8F03F8CF8CC1E3E73E0C33201E58C6F7F4F3E7E3003BBFC1";
    attribute INIT_20 of inst : label is "F800E003DE67B70301FC070C7C39007F81FB8446F03DE64CF7FC1F07E3983800";
    attribute INIT_21 of inst : label is "0F0071FF018FF8C01F0FF01F80067FC0383FFFF99E4CC0C9C0701F3EFFE001F1";
    attribute INIT_22 of inst : label is "1F800007E3FC0FFCF1E031C1F020C7FC3CFC707FFC007FFE70000E0FC387FFE1";
    attribute INIT_23 of inst : label is "FFFE00067FFFF80003C1FF8070000003FFFFFC00FFF003C03C01C10E71C3C71C";
    attribute INIT_24 of inst : label is "FC000007FFFE0003FF800FFFE0000FFFFE0700007FF1FFF803FF1FE380703C07";
    attribute INIT_25 of inst : label is "0003FFFFFFF10000060FFFF81C03F03F81FC0180047E00FFFE0FE0780E0001FF";
    attribute INIT_26 of inst : label is "01FFF0007FFE000FFFC001C7FFFFFF000F807C007C1FF007FFFFC0003FFF0000";
    attribute INIT_27 of inst : label is "FFE3DE0007FFFFFFF00183FFFEFC00000FFFFFF8000000FFFFF807FE0001FF80";
    attribute INIT_28 of inst : label is "DF00001FFFE007F807F801FE00FF801FF00FF001FFFFFC000607FFFFFFC0000F";
    attribute INIT_29 of inst : label is "000000003FFFF00000001FFFF0000F180003FFF800FFC1E003E703FFC780073F";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "D638DA1E4EF4CA4A15930237CD8D2442187B3F038FB4AAE7C1BC636D00E33ADE";
    attribute INIT_01 of inst : label is "B8D18C593C14EAA61566C15F61A97C7998836C268E713669CE386A3F438C7293";
    attribute INIT_02 of inst : label is "0E6DA6671A45B0F76946DD2D916398D88B61FCCF665CC8DE6C4932522E336F2C";
    attribute INIT_03 of inst : label is "66F9E961E9A0D93BACA650F39918E9198926DBE0EEE33325AE6608F3365A98CD";
    attribute INIT_04 of inst : label is "B9993B732CBFC59EE745F5753B3BB28F1DDB59BE322C6B1DAA27321DA4ADF559";
    attribute INIT_05 of inst : label is "24C9F8919BC0663472646736B4E6A54C732F18DCB9334D249E31B052669FA32F";
    attribute INIT_06 of inst : label is "F4F95287467683365C0CEF495A9875F613849472506C9DC659F674999B679269";
    attribute INIT_07 of inst : label is "40B28A6BE4D52E15F07F3EB86C4F393F10006C46E0FCB5431F97B612EE6EA744";
    attribute INIT_08 of inst : label is "6CAB5C5E2B1FBE6E7873B02E9207C416D2A614642926831CFBB560B5C27F38CA";
    attribute INIT_09 of inst : label is "DB64F336F9CDB6768A466588F4C582D81B3ECEAC544DB461686466950F46B674";
    attribute INIT_0A of inst : label is "92EEC308C5D866BBA2C3752B091AD29702A1DCD4555DF7049D644D11034B3534";
    attribute INIT_0B of inst : label is "80653FDD8BDD40CB1D13630CBE14A9E5C9AD32938ED7E9353DD64175936165CC";
    attribute INIT_0C of inst : label is "CF469A58EBA315F76258351716277C24A7CB41B2412CD2C9BD59F9075D23CA68";
    attribute INIT_0D of inst : label is "D4F2C70315F476776696497CB2D0524A2F30234BC89A90784F381BFFA5474D54";
    attribute INIT_0E of inst : label is "986DC92119962495EB76DDCA2A3288E22E684EFF53928C02AF378E24FBA74CF7";
    attribute INIT_0F of inst : label is "9CB3FCD3BF0FC893BD769726DE0CF6549161853B8F7BB8DA8CF2E385E3C595BF";
    attribute INIT_10 of inst : label is "5B039AB3113260E9FC2D2535E2FBEDD82E635D5B1A42EBAD1317EA4BB976D8D6";
    attribute INIT_11 of inst : label is "D84CE4156B5D46F735FF57BFB409E04CF253F8591914ECAF772C5887AD3295AB";
    attribute INIT_12 of inst : label is "3440255852764C84C974AB8424136ACD8FC191E4FF2104C3400DC2F9E49D602E";
    attribute INIT_13 of inst : label is "32AAC5BFCA8AAAD1637A3905B7818AD672C984C09D377B99FE27F8A99F75CB95";
    attribute INIT_14 of inst : label is "A40FC6F237F2BC79679F35087FA9BC4DBCEB58A0F33E0292D82AE58A334DF860";
    attribute INIT_15 of inst : label is "6A50FEDDFB4B8010E4E236ED83BC4AFCCAF380C3E310466D0875155ADB6DF636";
    attribute INIT_16 of inst : label is "342E5BEF8CF77794326ACBFE75FB4E380BC57E6DB7A97C5E0F165468CB2D5848";
    attribute INIT_17 of inst : label is "000DFB903B04CF4329529B3CACF90C8999303C7976003B985780C862A0D003B1";
    attribute INIT_18 of inst : label is "04E617FC8C0F33328216037E76F8200DEB0E60F03CBBCF91E007F28F8F8729D4";
    attribute INIT_19 of inst : label is "A17138E6770E018FCD8CF13326E7837523F06040073303E8F393F1E07D981C3C";
    attribute INIT_1A of inst : label is "DF9F6060733F2068070F20EE1E07CF80787D43719FF4FF81FC33BF9BE7DBF87F";
    attribute INIT_1B of inst : label is "9FF87184001E003031F982784C072013F3CF71FC00C7BFF1FF02660066E4E0C7";
    attribute INIT_1C of inst : label is "7F8F203C3C7F079FF0778FF80FC7C18033FC019F0DC0CFFE3C3F1F99CE78F67F";
    attribute INIT_1D of inst : label is "E063FC3FC3C000FF3E00001C0030FE7FE1F8303FE0007FFD9DF9F1C3EFF1C606";
    attribute INIT_1E of inst : label is "FF0000003FFFFEF010003FEFFFFC3C3FF7BF81FF1F807C1FE301C0001FF3077F";
    attribute INIT_1F of inst : label is "01FF01FF03F01FFF8F03F80F80FFFFE03E0C0C3FE1C7F8F80C0C07FF003FBFFF";
    attribute INIT_20 of inst : label is "F80000001F8070FC01FFFFFC03C1FFFF81F80047F03FFE4307FFFF00001FF800";
    attribute INIT_21 of inst : label is "0F0071FF018FF8001FFFF01F80007FC03FFFFFF87F8F00383F801F3FFFE001FF";
    attribute INIT_22 of inst : label is "00000007FFFC0FFCF1E00001FFDFC0003FFC007FFC007FFFF000000FC3FFFFE1";
    attribute INIT_23 of inst : label is "FFFE00067FFFF8000001FFFFF0000003FFFFFC00FFF003C03C01FFFE0E03F8FC";
    attribute INIT_24 of inst : label is "FC000007FFFE0003FF800FFFE0000FFFFE0700007FF1FFF803FF0003FFF00007";
    attribute INIT_25 of inst : label is "0003FFFFFFF10000060FFFF81C03F03F81FC0180047E00FFFE0FE0780E0001FF";
    attribute INIT_26 of inst : label is "01FFF0007FFE000FFFC001C7FFFFFF0000007FFFFC000007FFFFC0003FFF0000";
    attribute INIT_27 of inst : label is "FFE3DE0007FFFFFFF00183FFFEFC00000FFFFFF8000000FFFFF807FE0001FF80";
    attribute INIT_28 of inst : label is "DF00001FFFE007F807F801FE00FF801FF00FF001FFFFFC000607FFFFFFC0000F";
    attribute INIT_29 of inst : label is "000000003FFFF00000001FFFF0000F180003FFF800FFC1E003E703FFC780073F";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "3DC0E1063CBF038C147FE305F609C7062D570B3C0EAC7FE8009F838E4FE0FFEE";
    attribute INIT_01 of inst : label is "34BDBC8BCE8C37B86081C89FBAC71581E1971CDD0F962E187DC0760BFC0F388F";
    attribute INIT_02 of inst : label is "CDE39F781DF9704E1E42398E0CE5E0E1871868F231CAF101E36C3C609E0F1DCF";
    attribute INIT_03 of inst : label is "1E23C018AE39B8F37080600F81869C1E1961C7A6FB83CC1C60786070F1C720F1";
    attribute INIT_04 of inst : label is "2878F3E3CE8A67A4B16C7E21DF2A503CA9630873C71CB41B305F0E2460CDBA62";
    attribute INIT_05 of inst : label is "E397339DE30E1E5E20780F0E68DB3338C29AEA59823C671C70C1C3C1E18743CC";
    attribute INIT_06 of inst : label is "9C2F781CC078E6F1C78F3B399A1E62AE3687E83C631C79E79DCE19E04479C9F2";
    attribute INIT_07 of inst : label is "1771AC354BA76632AAD3CC2DE32BD71C1DF11D00E6592C0C2F8E617F550BE86F";
    attribute INIT_08 of inst : label is "7020E115E00AB5BA3DEB3CDF30B4060731E78B2A04E323D951F12BC08B5032BC";
    attribute INIT_09 of inst : label is "C71CC3C62D3C73B8E361E7AC7D87AB0A870EC28F9B7C72E59C5861B30ABA71EF";
    attribute INIT_0A of inst : label is "8E28EEE7F977068D64DDE7D8C553340672C6C095B56373E6CF78588D80C3C6FB";
    attribute INIT_0B of inst : label is "1578B36611A0E36656B0FBFDB15DC74CDE314EEAB719C70C3FDB9A938FE279CF";
    attribute INIT_0C of inst : label is "F30C79D98394D0C24C43E862561283BECBBF33DC61A3C78F94FF3E3741997619";
    attribute INIT_0D of inst : label is "195B023DA360B9D90E4071A171737B8C34F319AC22818F99996591A69C127D44";
    attribute INIT_0E of inst : label is "FA839FBF57E335A727B1C76C034672D5939A4C49408E3527A272DDC421BDA3C0";
    attribute INIT_0F of inst : label is "4A7283CCC17A2C19BCBC9A104E8F9190C8394CFA7B73971B8EDA4D4623FB88F1";
    attribute INIT_10 of inst : label is "93EB567344BDEA8DE7E43F3947280C824FEDC96B070146C24BF122B5377FE69C";
    attribute INIT_11 of inst : label is "C3DB57F2F3132F58DB88EFD0716FA00601A3F8E7401D8430D91EE09238967B69";
    attribute INIT_12 of inst : label is "683FE338640EDADD70D267F1680CA6310397B1F84030B9E0E8031E6FE3858018";
    attribute INIT_13 of inst : label is "EE66393FC7037334E3B9D983C75F715871F087A8DEBF887805C85F99F79BB0B6";
    attribute INIT_14 of inst : label is "9C083B0E38FD803E647038F0201BC1713FA6C720FC3F7C4E3833E671C820728B";
    attribute INIT_15 of inst : label is "E66701E380CC001B1DE9C0B1FF6C0CFC0C0180FE04F381E9F7F9F3CA138E2671";
    attribute INIT_16 of inst : label is "C7CE37F07700EFE7F18CC7FF8C07103FFC3B00618FC9803E000F9818F81E67CF";
    attribute INIT_17 of inst : label is "0001FC703F030F80E0CCDC3C63FEF137870FC3F9B800397867FFC79CC0300380";
    attribute INIT_18 of inst : label is "FC01E7FCFC0F00C301F1FC7E0707E003F3F1E0F000FC3F8000000CF07FFFE638";
    attribute INIT_19 of inst : label is "3E70F801F80FFFFFC070F1FCFE180086200FDFBFF83C00180FE3FFE001F81FFF";
    attribute INIT_1A of inst : label is "C0007FE07F3F1F8FFFFF1F0FFE000FFF87FCC381E00C0001FC3F801C1FF80780";
    attribute INIT_1B of inst : label is "1FF80E07FFFE00003FF87C7FF3FF1FE3FFCFF1FC0007BFFFFF0187FFE1F8FF3F";
    attribute INIT_1C of inst : label is "00703FC3FC00001FF07FFFF80FC001FFF00001E0FC3F0FFE3C3F1F860FFF0E00";
    attribute INIT_1D of inst : label is "E003FC3FC3C000FF3E00001FFFF0007FE0003FFFE0007FFD8001FFFFE001FFFE";
    attribute INIT_1E of inst : label is "FF0000003FFFFEF000003FEFFFFC003FFFFF80001FFFFC0003FFC0001FF007FF";
    attribute INIT_1F of inst : label is "01FF01FF03F01FFF8F03F80F80FFFFE03E0C003FFFC000FFFC0007FF003FBFFF";
    attribute INIT_20 of inst : label is "F80000001FFFF00001FFFFFC0001FFFF81F80047F03FFE4007FFFF00001FF800";
    attribute INIT_21 of inst : label is "0F0071FF018FF8001FFFF01F80007FC03FFFFFF8000FFFF800001F3FFFE001FF";
    attribute INIT_22 of inst : label is "00000007FFFC0FFCF1E00001FFFFC0003FFC007FFC007FFFF000000FC3FFFFE1";
    attribute INIT_23 of inst : label is "FFFE00067FFFF8000001FFFFF0000003FFFFFC00FFF003C03C01FFFE0003FFFC";
    attribute INIT_24 of inst : label is "FC000007FFFE0003FF800FFFE0000FFFFE0700007FF1FFF803FF0003FFF00007";
    attribute INIT_25 of inst : label is "0003FFFFFFF10000060FFFF81C03F03F81FC0180047E00FFFE0FE0780E0001FF";
    attribute INIT_26 of inst : label is "01FFF0007FFE000FFFC001C7FFFFFF0000007FFFFC000007FFFFC0003FFF0000";
    attribute INIT_27 of inst : label is "FFE3DE0007FFFFFFF00183FFFEFC00000FFFFFF8000000FFFFF807FE0001FF80";
    attribute INIT_28 of inst : label is "DF00001FFFE007F807F801FE00FF801FF00FF001FFFFFC000607FFFFFFC0000F";
    attribute INIT_29 of inst : label is "000000003FFFF00000001FFFF0000F180003FFF800FFC1E003E703FFC780073F";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "FD00FE9E03F003F043FA9E879C09F809FC10FFC00FB3FFEFFEA003F0181FFAFE";
    attribute INIT_01 of inst : label is "C000FC2FF01C0BBF879FC2BBEF10FF01FE0F03EA0FE81E07FE007EFF000FC180";
    attribute INIT_02 of inst : label is "03E07F401F5E5D418FAA078FE81F80FE2F07F0FD303AFE17E0BC3F81C1FF02AF";
    attribute INIT_03 of inst : label is "FE0EDF07CFC0780EB8AB80A07A817E1FE0E03FCB0103FC83E87F800FF03F00FE";
    attribute INIT_04 of inst : label is "27F80FC3F300977143FC059FEA7B479C63FC380CF883F01FC000FE03E8D3BF82";
    attribute INIT_05 of inst : label is "DE2F4875FC0DFE05FC7FE901E8C9C9077C1B8987883F8F03F901FC17E07F83F0";
    attribute INIT_06 of inst : label is "85AF2E53F87F01F03E0FC107211F859E22EE563F80FC0787E05E0700367E17FD";
    attribute INIT_07 of inst : label is "B4F057EAA85F2D50AAF9F09BE05C90FE1F2903E1B95723EFC181FF33D540C4FF";
    attribute INIT_08 of inst : label is "7F8813D2CB6BB9545C1F3F9FDBF998D48F07F63C941F03F6618E7A4FA5F6352F";
    attribute INIT_09 of inst : label is "C0F983F864FC0DBF06DFE59BDC074C0E7F033E8FE1BC0F9D40406070F34BF018";
    attribute INIT_0A of inst : label is "81C4E3A0019D075F1AC5F8983C63F29DAAF940FD88FF2B75B47F2A82FFF3F867";
    attribute INIT_0B of inst : label is "A67F93904277DB0BDAF013FC1F31B7234FC3BEC653E09F01C02BFC5F80BE7E49";
    attribute INIT_0C of inst : label is "FCF9F867D38DE7E1326BE46C340E213D0E810D5F849FC62F8D5F7FC63E2F2E07";
    attribute INIT_0D of inst : label is "1E63FE8190653FCB09C57E62F07023F093F006B01CF7801BEF43626F231ECC90";
    attribute INIT_0E of inst : label is "F9A06A3F300139389F703A700CD1FCCC2BF930309F9184C0DE4E417BE2C35FC0";
    attribute INIT_0F of inst : label is "39F3003EFE79E41D3C7D9C0F6E704FECEFB9DC060CA38FE670C22197E3D78105";
    attribute INIT_10 of inst : label is "1C0CCE0CC6C0198E081C3CC180180C43701E3B73007F81A06C0E1D83318080E2";
    attribute INIT_11 of inst : label is "C3C7980E031F1F9FE007DFE00E4F9FFDFFC3F880C0E3893FCB00809BC471FF12";
    attribute INIT_12 of inst : label is "B0001F0787FE39167FCE1FF1B00061FE001871FFC03F80000FFF1E0FE079FFF8";
    attribute INIT_13 of inst : label is "E1E1FE3FC003FC0C1C3819FFF8C0FF9F8FFF8798E0C007F803F06079F01F8077";
    attribute INIT_14 of inst : label is "83F003FE3FFF800067F03FFFE007FE7E3F9E3FDF003F803E07C3E7FFF81FFCF3";
    attribute INIT_15 of inst : label is "E187FFFF8030001C03E7FF3E00E3F0FC0FFF80FE07F00011FFFE0FC61C0FC60F";
    attribute INIT_16 of inst : label is "07F1F00007FFE007F00F3FFFFC00E03FFFFF00618009FFFE00001FF8F8007FCF";
    attribute INIT_17 of inst : label is "0001FFF03F000FFFE03F1FC3E00001C07F0000063FFFC70787FFC000FFF00380";
    attribute INIT_18 of inst : label is "FC0007FCFC0F0003FFF0007E07FFE00003FFE0F000FFFF80000000FFFFFFE000";
    attribute INIT_19 of inst : label is "3F8FF800000FFFFFC000F1FFFE000007DFFFC000003FFFF80003FFE001F81FFF";
    attribute INIT_1A of inst : label is "C0007FE07F3F000FFFFF000FFE000FFFFFFC3C01FFFC0001FC3F801FFFF80000";
    attribute INIT_1B of inst : label is "1FF80007FFFE00003FF8007FFFFF0003FFCFF1FC0007BFFFFF0007FFE000FFFF";
    attribute INIT_1C of inst : label is "00003FFFFC00001FF07FFFF80FC001FFF00001FFFC000FFE3C3F1F800FFFFE00";
    attribute INIT_1D of inst : label is "E003FC3FC3C000FF3E00001FFFF0007FE0003FFFE0007FFD8001FFFFE001FFFE";
    attribute INIT_1E of inst : label is "FF0000003FFFFEF000003FEFFFFC003FFFFF80001FFFFC0003FFC0001FF007FF";
    attribute INIT_1F of inst : label is "01FF01FF03F01FFF8F03F80F80FFFFE03E0C003FFFC000FFFC0007FF003FBFFF";
    attribute INIT_20 of inst : label is "F80000001FFFF00001FFFFFC0001FFFF81F80047F03FFE4007FFFF00001FF800";
    attribute INIT_21 of inst : label is "0F0071FF018FF8001FFFF01F80007FC03FFFFFF8000FFFF800001F3FFFE001FF";
    attribute INIT_22 of inst : label is "00000007FFFC0FFCF1E00001FFFFC0003FFC007FFC007FFFF000000FC3FFFFE1";
    attribute INIT_23 of inst : label is "FFFE00067FFFF8000001FFFFF0000003FFFFFC00FFF003C03C01FFFE0003FFFC";
    attribute INIT_24 of inst : label is "FC000007FFFE0003FF800FFFE0000FFFFE0700007FF1FFF803FF0003FFF00007";
    attribute INIT_25 of inst : label is "0003FFFFFFF10000060FFFF81C03F03F81FC0180047E00FFFE0FE0780E0001FF";
    attribute INIT_26 of inst : label is "01FFF0007FFE000FFFC001C7FFFFFF0000007FFFFC000007FFFFC0003FFF0000";
    attribute INIT_27 of inst : label is "FFE3DE0007FFFFFFF00183FFFEFC00000FFFFFF8000000FFFFF807FE0001FF80";
    attribute INIT_28 of inst : label is "DF00001FFFE007F807F801FE00FF801FF00FF001FFFFFC000607FFFFFFC0000F";
    attribute INIT_29 of inst : label is "000000003FFFF00000001FFFF0000F180003FFF800FFC1E003E703FFC780073F";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "FFFF0011FFF7FC0030047FEFB7F60008034FFF7FF00FFFCFFFBFFC00080004FE";
    attribute INIT_01 of inst : label is "008183FE0043FFC003403F74042FFFFE0010FFF3F00041FFFBFF83FF7FF0027F";
    attribute INIT_02 of inst : label is "081FFFFFE000603FD001FFB003FFBF0000FFEF002FFF00001FFDC0004000FFF0";
    attribute INIT_03 of inst : label is "01F452FFB00107FF0F5C0060047FFBE0011FFFF3FFFC017FFF8001000FFFBF00";
    attribute INIT_04 of inst : label is "0007FF7C017D0C6E8103EB7A04246203C68027FD017FF7E0004001FFFF36C000";
    attribute INIT_05 of inst : label is "40E087FE000401E3F78014FFFF3A04FE8044E5BFC3C004FFFDFE00001FFEFC00";
    attribute INIT_06 of inst : label is "7BF0E3CFEF80040FFEF004FE1DE00381C58D8F400203FFB800C1FE000B800FFE";
    attribute INIT_07 of inst : label is "0A0FE818E7E8E8CF24C200781F904FFBE0C4FFBFC0DCDFB0047FBF0436CE0820";
    attribute INIT_08 of inst : label is "8067E06E0CF6418FC3FDC0401C7E40C87FB80FE0F3FFBC0F808064379F8BCC30";
    attribute INIT_09 of inst : label is "3FFEFC001C03FEC001C01987E2F8F00600FC01300083FF027FBF9FF003860FFD";
    attribute INIT_0A of inst : label is "7FF71C6001E307C0FCC60047FE7C0E63CD00C0F27E80E3047980F67F001C0010";
    attribute INIT_0B of inst : label is "C78073F03C07C30C218FE3FC20F1871F90008101E40040FE000C00307FC38034";
    attribute INIT_0C of inst : label is "000407801C7C07FF018C1C600801C1C3F180FE60038039CF8260FFF90030E1FF";
    attribute INIT_0D of inst : label is "E07C01818F99C038F039801E0F8FBC00700FFF3FFF0F80180F7F03E03F1E33E7";
    attribute INIT_0E of inst : label is "079FF3C0F000C1C07F0FFC7FF03000C3CC0700001F9F8400FE7E3E7FE300C03F";
    attribute INIT_0F of inst : label is "F80C0000FF87E3E1C3FC600071FFC0030FC63C01F03C7FFE00C21E181C307E06";
    attribute INIT_10 of inst : label is "1FF03E0038FFF8700FFC3C01FFF80C3C7FFFF883007FFF9F8FFFFF80CE00FF01";
    attribute INIT_11 of inst : label is "C3C01FFE031F001FFFFFC00000707FFC0003F8FFC00071C038FF009C03F000FC";
    attribute INIT_12 of inst : label is "3FFFFF0007FE07E7803E000E3FFFE000001FF1FFC03F80000FFF1E0FE001FFF8";
    attribute INIT_13 of inst : label is "1FE0003FC003FFFC003819FFFFC0001FFFFF878700FFFFF800007FF9F01F8008";
    attribute INIT_14 of inst : label is "800003FE3FFF800067F03FFFE000007FC07E0000003FFFFE0003E7FFF80000FC";
    attribute INIT_15 of inst : label is "E007FFFF8000001FFFE0003FFFE000FC0FFF80FE07F00001FFFFFFC1E00FF9FF";
    attribute INIT_16 of inst : label is "07FFF00007FFE007F00FFFFFFC00003FFFFF00618009FFFE00001FF8F8007FCF";
    attribute INIT_17 of inst : label is "0001FFF03F000FFFE0001FFFE00001FFFF0000003FFFFF0007FFC000FFF00380";
    attribute INIT_18 of inst : label is "FC0007FCFC0F0003FFF0007E07FFE00003FFE0F000FFFF80000000FFFFFFE000";
    attribute INIT_19 of inst : label is "3FFFF800000FFFFFC000F1FFFE000007FFFFC000003FFFF80003FFE001F81FFF";
    attribute INIT_1A of inst : label is "C0007FE07F3F000FFFFF000FFE000FFFFFFC0001FFFC0001FC3F801FFFF80000";
    attribute INIT_1B of inst : label is "1FF80007FFFE00003FF8007FFFFF0003FFCFF1FC0007BFFFFF0007FFE000FFFF";
    attribute INIT_1C of inst : label is "00003FFFFC00001FF07FFFF80FC001FFF00001FFFC000FFE3C3F1F800FFFFE00";
    attribute INIT_1D of inst : label is "E003FC3FC3C000FF3E00001FFFF0007FE0003FFFE0007FFD8001FFFFE001FFFE";
    attribute INIT_1E of inst : label is "FF0000003FFFFEF000003FEFFFFC003FFFFF80001FFFFC0003FFC0001FF007FF";
    attribute INIT_1F of inst : label is "01FF01FF03F01FFF8F03F80F80FFFFE03E0C003FFFC000FFFC0007FF003FBFFF";
    attribute INIT_20 of inst : label is "F80000001FFFF00001FFFFFC0001FFFF81F80047F03FFE4007FFFF00001FF800";
    attribute INIT_21 of inst : label is "0F0071FF018FF8001FFFF01F80007FC03FFFFFF8000FFFF800001F3FFFE001FF";
    attribute INIT_22 of inst : label is "00000007FFFC0FFCF1E00001FFFFC0003FFC007FFC007FFFF000000FC3FFFFE1";
    attribute INIT_23 of inst : label is "FFFE00067FFFF8000001FFFFF0000003FFFFFC00FFF003C03C01FFFE0003FFFC";
    attribute INIT_24 of inst : label is "FC000007FFFE0003FF800FFFE0000FFFFE0700007FF1FFF803FF0003FFF00007";
    attribute INIT_25 of inst : label is "0003FFFFFFF10000060FFFF81C03F03F81FC0180047E00FFFE0FE0780E0001FF";
    attribute INIT_26 of inst : label is "01FFF0007FFE000FFFC001C7FFFFFF0000007FFFFC000007FFFFC0003FFF0000";
    attribute INIT_27 of inst : label is "FFE3DE0007FFFFFFF00183FFFEFC00000FFFFFF8000000FFFFF807FE0001FF80";
    attribute INIT_28 of inst : label is "DF00001FFFE007F807F801FE00FF801FF00FF001FFFFFC000607FFFFFFC0000F";
    attribute INIT_29 of inst : label is "000000003FFFF00000001FFFF0000F180003FFF800FFC1E003E703FFC780073F";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "FE00000FFFF800000FFFFF1FC8000007FFBFFF80001FFFF00040000007FFFF01";
    attribute INIT_01 of inst : label is "007E7FFC003FFF00003FFFF8181FFE00000FFFFC00003FFFFC0001FF800001FF";
    attribute INIT_02 of inst : label is "07FFFF80003F80FFE007FFC007FFC0001FFFF0001FFC000FFFFE00003FFFFFC0";
    attribute INIT_03 of inst : label is "FFF821FFC000FFFFF000001FFFFFFC0000FFFFFC000000FFF00000FFFFFFC000";
    attribute INIT_04 of inst : label is "1FFFFF8000FE039F00FFF0FC001F81FFFF001FFE00FFF800003FFFFFF00F0001";
    attribute INIT_05 of inst : label is "3F1FFFF80003FFFFF80003FFF00403FF003F1E7FFC0003FFFE00000FFFFF0000";
    attribute INIT_06 of inst : label is "FFC01C3FF00003FFFF0003FFFE00007FF873FF8001FFFFC0003FFFFFFC000000";
    attribute INIT_07 of inst : label is "01FFF0071FF0103FDF3C0007FFE03FFC0003FFC00023FFC003FFC0F80831F01F";
    attribute INIT_08 of inst : label is "001FFF81F001FE003FFE003FE0003F3FFFC0001F0FFFC000007F9FF87FFC03C0";
    attribute INIT_09 of inst : label is "FFFF000003FFFF00003FFE7FFF000001FFFFFFC0007FFFFF8000000FFC01FFFE";
    attribute INIT_0A of inst : label is "FFF8001FFE00F83FFF38003FFF8001FFF0003F0FFF001CFBFE0001FFFFE0000F";
    attribute INIT_0B of inst : label is "F8000C0FFFF83CF0007FFC03C00E78FFE0007FFFF8003FFFFFF0000FFFFC0003";
    attribute INIT_0C of inst : label is "0003FFFFE003F800FFF0039FFFFFFE00007FFF80007FFFF07F800000FFC01FFF";
    attribute INIT_0D of inst : label is "FF80007E7FFE0007FFFE0001FFFFC0000FFFFFC000007FE7F080FC1FC0E1FFF8";
    attribute INIT_0E of inst : label is "007FFC000FFFFE0000FFFF80000FFF3FF000FFFFE0607BFF0181FF801C003FFF";
    attribute INIT_0F of inst : label is "07FFFFFF00001FFE0003FFFF80003FFFF00003FFFFC00001FF3DFFE0000FFFF8";
    attribute INIT_10 of inst : label is "E00001FFFF0007FFF003C3FE0007F3FF800007FCFF80007FF000007FFFFF0000";
    attribute INIT_11 of inst : label is "3C3FE001FCE0FFE000003FFFFF800003FFFC07003FFFFE0007FFFF60000FFFFF";
    attribute INIT_12 of inst : label is "C00000FFF801FFF80001FFFFC0001FFFFFE00E003FC07FFFF000E1F01FFE0007";
    attribute INIT_13 of inst : label is "001FFFC03FFC0003FFC7E600003FFFE00000787FFF000007FFFF80060FE07FFF";
    attribute INIT_14 of inst : label is "7FFFFC01C0007FFF980FC0001FFFFF800001FFFFFFC00001FFFC180007FFFF00";
    attribute INIT_15 of inst : label is "1FF800007FFFFFE0001FFFC0001FFF03F0007F01F80FFFFE0000003FFFF00000";
    attribute INIT_16 of inst : label is "F8000FFFF8001FF80FF0000003FFFFC00000FF9E7FF60001FFFFE00707FF8030";
    attribute INIT_17 of inst : label is "FFFE000FC0FFF0001FFFE0001FFFFE0000FFFFFFC00000FFF8003FFF000FFC7F";
    attribute INIT_18 of inst : label is "03FFF80303F0FFFC000FFF81F8001FFFFC001F0FFF00007FFFFFFF0000001FFF";
    attribute INIT_19 of inst : label is "C00007FFFFF000003FFF0E0001FFFFF800003FFFFFC00007FFFC001FFE07E000";
    attribute INIT_1A of inst : label is "3FFF801F80C0FFF00000FFF001FFF0000003FFFE0003FFFE03C07FE00007FFFF";
    attribute INIT_1B of inst : label is "E007FFF80001FFFFC007FF800000FFFC00300E03FFF8400000FFF8001FFF0000";
    attribute INIT_1C of inst : label is "FFFFC00003FFFFE00F800007F03FFE000FFFFE0003FFF001C3C0E07FF00001FF";
    attribute INIT_1D of inst : label is "1FFC03C03C3FFF00C1FFFFE0000FFF801FFFC0001FFF80027FFE00001FFE0001";
    attribute INIT_1E of inst : label is "00FFFFFFC000010FFFFFC0100003FFC000007FFFE00003FFFC003FFFE00FF800";
    attribute INIT_1F of inst : label is "FE00FE00FC0FE00070FC07F07F00001FC1F3FFC0003FFF0003FFF800FFC04000";
    attribute INIT_20 of inst : label is "07FFFFFFE0000FFFFE000003FFFE00007E07FFB80FC001BFF80000FFFFE007FF";
    attribute INIT_21 of inst : label is "F0FF8E00FE7007FFE0000FE07FFF803FC0000007FFF00007FFFFE0C0001FFE00";
    attribute INIT_22 of inst : label is "FFFFFFF80003F0030E1FFFFE00003FFFC003FF8003FF80000FFFFFF03C00001E";
    attribute INIT_23 of inst : label is "0001FFF9800007FFFFFE00000FFFFFFC000003FF000FFC3FC3FE0001FFFC0003";
    attribute INIT_24 of inst : label is "03FFFFF80001FFFC007FF0001FFFF00001F8FFFF800E0007FC00FFFC000FFFF8";
    attribute INIT_25 of inst : label is "FFFC0000000EFFFFF9F00007E3FC0FC07E03FE7FFB81FF0001F01F87F1FFFE00";
    attribute INIT_26 of inst : label is "FE000FFF8001FFF0003FFE38000000FFFFFF800003FFFFF800003FFFC000FFFF";
    attribute INIT_27 of inst : label is "001C21FFF80000000FFE7C000103FFFFF0000007FFFFFF000007F801FFFE007F";
    attribute INIT_28 of inst : label is "20FFFFE0001FF807F807FE01FF007FE00FF00FFE000003FFF9F80000003FFFF0";
    attribute INIT_29 of inst : label is "FFFFFFFFC0000FFFFFFFE0000FFFF0E7FFFC0007FF003E1FFC18FC00387FF8C0";
    attribute INIT_2A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_31 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_32 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
