-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "44A212717677EC30C1A49428B1054B47FF8451F4A891B426532EDB1795E00799";
    attribute INIT_01 of inst : label is "98AC7B4EA7E89B7353567E0A86089A3C4A16806BC3C60C1E3C70F08FFF56B915";
    attribute INIT_02 of inst : label is "F554F2411434700F4146CC6416A712CC92F37E8E88000EB3CC51C54731431E05";
    attribute INIT_03 of inst : label is "9A851C6633F52D1389865F9E8BB3EAE299A261D2A418497E25C51677EDE93674";
    attribute INIT_04 of inst : label is "B001B3F3B315710D1A5D87EC4E92EC475008AA69C43DDD75B7CB220108EABCE2";
    attribute INIT_05 of inst : label is "D54C0E8198A8D3FB9C5000B5002FCED32A1DDF276CA63A8A859472776B80A100";
    attribute INIT_06 of inst : label is "C11A11614C15CFCFA6F3ECFF3F84C41682A00928C5AE148394219CB975E79194";
    attribute INIT_07 of inst : label is "B9C8C9C85D91BB7549778E2825DCCDC2DE9193EFB27A7E4F1AB4782DECC83390";
    attribute INIT_08 of inst : label is "01F218B13AD806D84DAF34935CB500AA8877BDF783EABC3870101C84D7885920";
    attribute INIT_09 of inst : label is "DE50E10C6215B3E15F52158D18D14200BB23EAD2447CBCF5ED90A8666632CC3D";
    attribute INIT_0A of inst : label is "2BA01737A2C7959598BDB93D12B30B93F51ABEAB5DD6F722FEB11CB86B422234";
    attribute INIT_0B of inst : label is "D00022D25B216AA256E2A0D6D7052050D4AD9DD0F9FD234EAEB0A1547BD7740A";
    attribute INIT_0C of inst : label is "61A97A5A001114315D4C498A31112B5956CDFD985E6D2AA222974D65C541AD5A";
    attribute INIT_0D of inst : label is "03FA2C45528A45EC1EC10806916BA53A7F644D78CC6A83BAAB28A077BD8053A0";
    attribute INIT_0E of inst : label is "6DF7E9730303135445F31355664B8EEC16631895C57D22A5DCE869703D095F59";
    attribute INIT_0F of inst : label is "223BFA9CD6C9008055561578768F63BA574676214DE3CF73DCDA5888FA2774E9";
    attribute INIT_10 of inst : label is "E064E51C0CBF4CC4735988EA713A98E62074080A00907DF71ADD296810128811";
    attribute INIT_11 of inst : label is "BBE62703E3FED383BC14CFFB8857EED266DB78D3E69F36F9B9305DDABE33D9CD";
    attribute INIT_12 of inst : label is "29448FD6EEE94E9674FFC9AFFF5C2E27DFDFC48F32FFFD3F5959DEBA79DC4525";
    attribute INIT_13 of inst : label is "10024CF020397CDF9BABE055B390E88A49E71963B20F84011EFF9991EC77237A";
    attribute INIT_14 of inst : label is "235EB5758FDFB2A3F9B65F85FFB31FFF72EB89008352D5A662159D34AAC3BBBF";
    attribute INIT_15 of inst : label is "DDD7775C2A0982510108822DA5EB07B95552AA0B895555A9B54769E3B41FC906";
    attribute INIT_16 of inst : label is "DD75DDDD6AFB5775DD556D55D5555A94C55557606AFBABED7F5D742A097DDF75";
    attribute INIT_17 of inst : label is "F907CFF1CCADCB2D12AAA6D49AA752ABAAAAD29ACD54A1D2D564DF5D5F7F5555";
    attribute INIT_18 of inst : label is "A00007400937C060EAA5995F69BA2F2830A20AB5C63690E28A4C72C0E4B86A4D";
    attribute INIT_19 of inst : label is "D6EAEFEE7C045447BBAFAFAE77398A5B1C75386BF1BEAB0A950680E8A6CDEDAB";
    attribute INIT_1A of inst : label is "4141415850520405D2CDB0B32C6C2C857212003C1F0F83C3EB737AF4C441106E";
    attribute INIT_1B of inst : label is "000451082A00E452A2ACA8A8A8AA90651942C0B43414250514B8BB262E2E2EA1";
    attribute INIT_1C of inst : label is "31115F5FBFDFDE92FE37FFB7DE973F9EAEA577F0000C000FFC0FF00F00000000";
    attribute INIT_1D of inst : label is "24A70904AE3CC820046347290838045021C200A1E289199C0A1BAB6693754843";
    attribute INIT_1E of inst : label is "A9477CEFBA79DD15F457BB2B2964E48FFD59FB9CE7B0EC170808F7CF9FD06109";
    attribute INIT_1F of inst : label is "902546F6D6995CE591856337C5BFEC60CFECF4410F67F9C2DAFD18039DAA858A";
    attribute INIT_20 of inst : label is "60407FD962050003F310081036CB9A4CD6CDB7197094851950A398AB84DE2CC9";
    attribute INIT_21 of inst : label is "D8220678806409E2211AF41E003880F47FEC8A208FFA08391628840073FC5214";
    attribute INIT_22 of inst : label is "0AA7121D98044C99ECE67032720D065FA793B3A62FD5BFDFF70209C8B1401085";
    attribute INIT_23 of inst : label is "DDDD5DD7D3939287F87E3F1AF8FF7E91FBE05B74D11A64B3C45848DECE207710";
    attribute INIT_24 of inst : label is "4224A00004A5080000000000000003FFFFFFFFFFFFF9F0081A0827007FFFFFFF";
    attribute INIT_25 of inst : label is "006110A00919001020108C820001460C09320800103400004C10209144C68624";
    attribute INIT_26 of inst : label is "0108C52051091050420C000008110000B99018002C200A210640520044805478";
    attribute INIT_27 of inst : label is "7F7C414802884EE24300F0509680DB0300000000000000000000000000002538";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "B66727F2484910C3080026E47260A6880412301B76E7261022932C80221807A8";
    attribute INIT_01 of inst : label is "51C0FE507486738A7469401D5479D6025369CFB52A55AA52A5469E60007104A8";
    attribute INIT_02 of inst : label is "01F2801A71E3B0011A1C00C0346060830080555110B9426028E3F2F8A38E448A";
    attribute INIT_03 of inst : label is "01B639A4A0729F7635D404813242860D2BCC82499399028AC30348090924A410";
    attribute INIT_04 of inst : label is "65BDF88A40621D9A28C4D0A6B405A6348AC160160EF1B2D848822EECBB6D84BF";
    attribute INIT_05 of inst : label is "BE9352AA03114E04008F966869D65FA475A045473D50E4B4581DB5B8842C3596";
    attribute INIT_06 of inst : label is "8A2363658C9693089900500823F2D98C1F92C119D8A4CADE66B66000CE4B652F";
    attribute INIT_07 of inst : label is "6103201AA5060C069689155116A04BCC04813DF130C483B3BF5A9FD140C9440A";
    attribute INIT_08 of inst : label is "6C00DB43A32088A3B603896C6006983D1E87B40B155000AB33CCED1919359204";
    attribute INIT_09 of inst : label is "60CB64B99B5D468A82AD6E76A3066C59B85AC50B398EFA8B2486458CA0519085";
    attribute INIT_0A of inst : label is "F4CDEA8134A60A5A21440A31A3541448A23952586125108D8806602323BBCC4B";
    attribute INIT_0B of inst : label is "2673CD88AEC69700A98D042918D2B4FFEFB0042D13FCC4921325939994A0022E";
    attribute INIT_0C of inst : label is "ACB8C484DA2E60C2A435069427E6B4822A0319FC30A244CCCB1C921B1A0852E6";
    attribute INIT_0D of inst : label is "1CD39D88A1148A71E30E3121268E49E4881E8A4D5994CD485271C7B9454DE33D";
    attribute INIT_0E of inst : label is "800C12946A642DA9A66D65A980A2E515451D616E3E825F5A10039209C633A636";
    attribute INIT_0F of inst : label is "10A2046450026909A77D27ACA0C6905B6AD80C6CC30518CE314486F6D4CFC905";
    attribute INIT_10 of inst : label is "D2AE2CB3509492994A25128D46A152945D4395A73B4B0005E090BCEAA24B9E81";
    attribute INIT_11 of inst : label is "20178668EC0023DFDEFB1802658C422D09459300804402202CBDE4111FBEDFD9";
    attribute INIT_12 of inst : label is "6A9913B92AA9020AC908650BD4AD4A14966E22DF24AA80900405DDC48623985A";
    attribute INIT_13 of inst : label is "324EE32951A1050C82390B2020352B911FAB48A6A0DFB69772F20CB998AC05C8";
    attribute INIT_14 of inst : label is "452006C0106003468A01805A0200A00600112523ED2926000CE202491D144101";
    attribute INIT_15 of inst : label is "5D5D7577FD5755FBEBD5DD70F8BB5375999B315D2DE99A33BB6E338FDA711B28";
    attribute INIT_16 of inst : label is "FDD75557D07FF55D57FFD2F77FFFF2FE4FFFDD74507F41FFFD577FFD5755D577";
    attribute INIT_17 of inst : label is "78F7D7FEA5315C39C3CCD4A7A33C6B3273239CC35666C463664E13FFFFFFFFFF";
    attribute INIT_18 of inst : label is "B0000560F906C1E099C2BA0E3E05B6011C4014F6067E3D01CE206AC04E684F3F";
    attribute INIT_19 of inst : label is "54150550D7FAFFAFAFAAFAAF7F0D047B20F341EC3D19B5CD27B0401482EBFD87";
    attribute INIT_1A of inst : label is "20282030080C131260791E1E6767A78636160803FF0FFC000C0BA103C5014410";
    attribute INIT_1B of inst : label is "557540000001108052589595949704C4240D53109090C030390D0E4B43C303C8";
    attribute INIT_1C of inst : label is "582CE1144221555A30A02C08E3A18D47C672DFFAAA9CAA9FFEBFF2BF155FD855";
    attribute INIT_1D of inst : label is "DB56FECE61ABB64A3E489095AF36A7EF35BF35DAAEDEC5AE777235516E1CE5EB";
    attribute INIT_1E of inst : label is "722D9F94D797637F9DA8C8FE72093B80002000238CE42AA6F3290C081069DAD6";
    attribute INIT_1F of inst : label is "274BD09B783268C7241F98DA62039B0D930332AEA98062B5800CF7FCF6755A7F";
    attribute INIT_20 of inst : label is "1C2F98334DB1BDECCB5B67FACDB26D926DA2D75275282A439F3F8413A15F08DC";
    attribute INIT_21 of inst : label is "4F77791277A2D449DEA4AE85DF577D62D555559AD461F7C4A1456FDA0DC3AFE9";
    attribute INIT_22 of inst : label is "F9C7857A8B56835F6FEDE957165AA84A486056C9CC39A1146CBDF2250A2DBFE8";
    attribute INIT_23 of inst : label is "16340A02A802A8075AD6D68E89DF810502E4FFF7FBBFFF50FEFFFE1203F7ABFB";
    attribute INIT_24 of inst : label is "005103F2C010640000000000000003FFFFFFFFFFF552B55AB98C97D579143616";
    attribute INIT_25 of inst : label is "1880480D40405008010400510C80A10000002450200980A000400C42B029098A";
    attribute INIT_26 of inst : label is "40C5081F00008D0218608080100C69C24048E4008302000A010000202240A000";
    attribute INIT_27 of inst : label is "CC0FFCE77BEDB317B4AB5D2BCB696A7500000000000000000000000004000280";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "268B47F02222241042A024A261602247F80118C64CC35C0AF83C920630640784";
    attribute INIT_01 of inst : label is "48CC7F58B2E8BBC917092F0F9200FC747A48C424B93264C9972A5204051AA565";
    attribute INIT_02 of inst : label is "06544B501120B805D054006574303445AA50299998E947982461ED6C9181778B";
    attribute INIT_03 of inst : label is "0087B54399008103AD035AD5A95AA3EBF1EA30C08090404425440202A465123E";
    attribute INIT_04 of inst : label is "A94828199177B9977888F006B0848610C2A27A1226BD69EDF3D940042273B443";
    attribute INIT_05 of inst : label is "F7D5542A0999C45280DD1CFE7B6C5037BEAC4B7455438EA555ED3B84C5A02404";
    attribute INIT_06 of inst : label is "4B0945498914E4618BD4BD7187109002C2A40183900443D134A4D42A7B7DB5BC";
    attribute INIT_07 of inst : label is "388A129ADA45B536D62BD46A16D454260498B7FD32A6C0FF3BFAB169CEA96132";
    attribute INIT_08 of inst : label is "4A089271839C8CF2DF6FCDBE5414942F8AAFF0062B59B55E2199BB8F8FD8FA21";
    attribute INIT_09 of inst : label is "F0F3CB3553D5E552D15AD290B2B568120AF041501D7E068CA004012A6834D57A";
    attribute INIT_0A of inst : label is "7E48FE113EF13C9F0B508B89B3F13532531E640B86B2BFEAA7F544720ED1EA8D";
    attribute INIT_0B of inst : label is "5C51EBF1B9F369BCB75EB7368D19CF2148B083F553AB6ED9F9F772DDDE722666";
    attribute INIT_0C of inst : label is "293B36CA8A2F562B78F9C737E2F5BB5E5A00D934CEA36FEE6FD2DD7CBD6E6D38";
    attribute INIT_0D of inst : label is "96F31958F336DB3DB7DB9825B4E96C96F166CBEFD9DEE9E66FD166FDE4CCF884";
    attribute INIT_0E of inst : label is "A41FFEB54D6F76DDE7373EDDC28D4DF81A5E7BB9F3DB7B78B812DB69679BD7CF";
    attribute INIT_0F of inst : label is "71915E6118F349DD311EA1AC22C65052775002A8D8EB5AD6B546DA3C3E6F2D85";
    attribute INIT_10 of inst : label is "36EB29A85D8ADA4D29349A5F2793CA53E125AD694A5225EEA2552C42A4908C02";
    attribute INIT_11 of inst : label is "15C0815A08A091D5CEA91FF3CD954A6338CFD291088844423D38EC033F946BD4";
    attribute INIT_12 of inst : label is "03C03BB95555A306AD97656BCAE168525CBE643A14555106D8DDFE26FA8FD509";
    attribute INIT_13 of inst : label is "26CEB1D975187743A1C3C9250435D28C9FD42F61489126814CEC017984620328";
    attribute INIT_14 of inst : label is "01FAD32DA8689BE0AB508F8AFAD0AF9510F60F79472BF3D076B81B6DCFD57909";
    attribute INIT_15 of inst : label is "5FF57FDDDDDD77551475F570A0BEF9DE1E1C3D9E318E1CC2A84BCD037B1D1B06";
    attribute INIT_16 of inst : label is "DF7DFFFD453F7FFFFFD7D0FDFFFFF0D597FD778B853F14FDDDDFDDDDDDF5FD7D";
    attribute INIT_17 of inst : label is "8407D1FF05CE5FC1FC0F04B823C58BC243CC9F0BF87908787806FFDD7F7FDD5D";
    attribute INIT_18 of inst : label is "C00000500930207E4C94F1D9CC1E70CA75D2BF79272F7693B7C210E02D601689";
    attribute INIT_19 of inst : label is "54200D405600D40455AA80052BEADD1F923F247386C24B135B4F40794CE51E58";
    attribute INIT_1A of inst : label is "00000808020181811407020120E0E040C202090000F00003E9E2DFF8C40B2000";
    attribute INIT_1B of inst : label is "083100001010016062649A9B99988324D032CCB3333328C8C613114444044428";
    attribute INIT_1C of inst : label is "784A3F5998CC18C90EB21318030398C8E231CFFE101CAA9FFC1FF01F42222520";
    attribute INIT_1D of inst : label is "D6F9BEB2C71685928F91A3CF734CA9FB676F45D10D1E8E19B583C2B34839EE2C";
    attribute INIT_1E of inst : label is "3AB42D0F9DC4C42AE5AF2C553A10FA07B900F40A10284A65CEE23031E3D9B7BC";
    attribute INIT_1F of inst : label is "05B89418E345600648ACD1474395A2C6A45A5675C64889270C55D19BE1ED2955";
    attribute INIT_20 of inst : label is "03083B9A6B042201D842081096DC82E416CB21D2152C2B4650208E20A10F0658";
    attribute INIT_21 of inst : label is "086A120C05202830144A1C02148852052ADD8674D8892A38408A42B40A40230D";
    attribute INIT_22 of inst : label is "00B38F258A96E54A35EA1B7594542EC56C31A3283A172C72160A98C204501AD0";
    attribute INIT_23 of inst : label is "FEA8200A2220888FCE73A8DA6BB78184F9258926244B163141482DB206A81554";
    attribute INIT_24 of inst : label is "840A4001084A120020000000000003FFFFFFFFFFFF0E7F087BA692AAFFABFE89";
    attribute INIT_25 of inst : label is "20162000A082A0A1004902042000004202400308884009060221002401001041";
    attribute INIT_26 of inst : label is "04002040001062A5809108102522802400250210105C00003001040108080087";
    attribute INIT_27 of inst : label is "FADE49294AC1088F0528875A54BA865400000000000000000000000000804840";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "6240320B63C3A49A4AA2202D73E0226A8251100C4CE38462898C9B0611400780";
    attribute INIT_01 of inst : label is "9CF603BB37319CD3918B72CDA784CD939C8BE4998B060C583560DAC50510252C";
    attribute INIT_02 of inst : label is "2342D6405144B0034044036758A0B0E582F02CCCCBC446B04E7854FDB9E11A2F";
    attribute INIT_03 of inst : label is "43316CE63504B26C9896CC949B952EA8B662A89A84E940C0B03323A3AE54B7B4";
    attribute INIT_04 of inst : label is "231C000B1355A859180D842C00A52CA142006A0456695FFEDAFB6AE5A3689004";
    attribute INIT_05 of inst : label is "4ED6D6029888C869A2AD3DCE33684F96F728C26B4F1202191925B18361000D20";
    attribute INIT_06 of inst : label is "FB087164FCC7265932F0AC5D6456CC074A1002B758435D9BB1130D78232C9CD0";
    attribute INIT_07 of inst : label is "10FB52481F82966EC0327848070D47CE8471921B0EF2FED9EF7C234CE5D7619A";
    attribute INIT_08 of inst : label is "23F859AEA8CBDE38DB2465B7CD58195DACBC55F5CACC94B8F2A8BDADC4D8CCE5";
    attribute INIT_09 of inst : label is "BE55E14CD7587166C5AF7BDEBAF74E83801806400CD8C035E382046743A4553F";
    attribute INIT_0A of inst : label is "670ECF3477756FFB3C5DA72FF76745DF5378808A1597B52734937D19D0556665";
    attribute INIT_0B of inst : label is "95DD6656B9627898A77C9627C77AD6BDEF79A53979FD665D8D923AC4731BAAB7";
    attribute INIT_0C of inst : label is "095562D3ABEB327C4B5E5B97E2B3A3CB0E518B9D5861722364A65F2EF92C4F1C";
    attribute INIT_0D of inst : label is "D73755EAB5538B8DBCBBD97CB7F32EB2F3FEE329CAD62F3209857EE7320DDAAC";
    attribute INIT_0E of inst : label is "ED1E98B9C3F212C4599212C4760B4C8A165EF5BA62D17760CE50CB2B7159194B";
    attribute INIT_0F of inst : label is "603B927018620F8CD51C05F97446000B460E86C8A9895AD6B5C2CAB8B36065D7";
    attribute INIT_10 of inst : label is "32C1A3A85A8A5CD47B59A8E37938DAE6207694AD294A35BA32E524602424CC09";
    attribute INIT_11 of inst : label is "3D76B66206A0B850606C4859DDB541CCD1C2D1B109884C409D03DC977F61A105";
    attribute INIT_12 of inst : label is "E8151DF47FF8E58465D5E6A56A7C68574C9F600FB85553024E4E72C2C8A8CD43";
    attribute INIT_13 of inst : label is "AF6C159D6C185C4A618369B5B59879BB0DC6454FF0402B3605054DD68D874D7C";
    attribute INIT_14 of inst : label is "A64C912488C83F61BD9528F28E9508D23453D6BD56ACB145C6357165BD91892B";
    attribute INIT_15 of inst : label is "5FFD7FFC002308EAAAF5E82A0895ABA81FE03E103E0FE0FC120E6543EB3BCD66";
    attribute INIT_16 of inst : label is "BBFFFFFF8010FFFFFFFBC2FFFFFFFF7A8FFFBFAA801000415577F40023F5FD7F";
    attribute INIT_17 of inst : label is "03330CFF500F5FFE270FFB42C309F3FD83F01BF403800300784E1EFBFAFEFFFF";
    attribute INIT_18 of inst : label is "A008042C071246622890101809341C0430511070A42EF451AE0A01C00C500E4D";
    attribute INIT_19 of inst : label is "097550950355095000DDDDD08318051A0A331461E0660300931100D280610D20";
    attribute INIT_1A of inst : label is "90908080202489880043121064E4A4110404000000000003E95D5FF6D95CF555";
    attribute INIT_1B of inst : label is "DDE000000404000042409190909002148020C8723232188881111084C4844408";
    attribute INIT_1C of inst : label is "3047116DD2E9AF5C285B5ED8A1CEFCFF5B9F9FFEBABE003FFEBFFBFF37FFF8F5";
    attribute INIT_1D of inst : label is "DCE912E79E9C3799898D9FE6B5C8DA95C644E44FE5126E7B19E55EBB23B9DEEC";
    attribute INIT_1E of inst : label is "5620819FC990E6A2788FBC45D601398AC68800808220121BA7845A34E9FCAF5B";
    attribute INIT_1F of inst : label is "33AE9428A112A00407A84FC743D0195D1179167F9F602F9B2D45A75E416D3925";
    attribute INIT_20 of inst : label is "8349785A2B646AD3D85AC854B6D8A6C532CB705105060922D1220C2621468E00";
    attribute INIT_21 of inst : label is "99045C180560B0601568A48614D8534D2A9D86F1D889096050D8461420202124";
    attribute INIT_22 of inst : label is "52B1072500DEC430D0829960D1542D452E300A648D11E2D29302580286C31850";
    attribute INIT_23 of inst : label is "CD98AAA888880007FFC2208820B7C0C18102A5AF202F9720082C3E844044C022";
    attribute INIT_24 of inst : label is "43A4A7F00321480000000000000003FFFFFFFFFFFF307F307D55582AFAF998CC";
    attribute INIT_25 of inst : label is "020116D2040108120022800A00280024CC08000514203640100C00090080A024";
    attribute INIT_26 of inst : label is "800A003F1A0500500000000800101200109011420C009C200400598090000060";
    attribute INIT_27 of inst : label is "9399D69CA73CFDF0D7A4ADFD757EA69500000000000000000000000000002104";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "E8CC700258593AE388C28B446B62B42AA95BA859767C4B5822B80009A8280781";
    attribute INIT_01 of inst : label is "0DCE8058526602C92B28265DE385DCB6592AEC108952240814205244A52B84F1";
    attribute INIT_02 of inst : label is "965684000042B008829041010844812408B2A9999CC6A50226EA4D6C1BAC064B";
    attribute INIT_03 of inst : label is "039324744102112D8C14A6070CD325209562A2C916959380767728293345A928";
    attribute INIT_04 of inst : label is "57BF659C17FFF063BA4FE23E45033E440A85541C1640804900124004A26D030B";
    attribute INIT_05 of inst : label is "86C407207DDDDA499B9C302CA5764D36B60BDB65107240921801B41832081C92";
    attribute INIT_06 of inst : label is "4BA0664CA99252499432A15D36128908D2B007911C26481CE2144C99636DBDB1";
    attribute INIT_07 of inst : label is "B210C35C6A94C5E6C8A4DBF2074C981598AB021E2456C1986370A4F18C8B743A";
    attribute INIT_08 of inst : label is "4E1A9111819BACB8736C64E64C845C2D9028580A9559B460673339EDCDDAD849";
    attribute INIT_09 of inst : label is "B001C404574D6552C14A4214B0A10C49C81D465B6C5042827934654DA6D7849A";
    attribute INIT_0A of inst : label is "662CCCF336E0AD5B06579B01BB70E5205B3910D4C468A96325B10CC980556224";
    attribute INIT_0B of inst : label is "E91462C6B47B81DCB93F56380C3084294AB792304FA86C4A1A3066CCD6301324";
    attribute INIT_0C of inst : label is "2B33827D2C8B1699991AEB5608B12C227B4A1136E1693667759848887EAC7031";
    attribute INIT_0D of inst : label is "F667198CB916AB1BB5BB5BA9B04C26C2501ECB7980D62D6633897EED66DFD015";
    attribute INIT_0E of inst : label is "9C949CAB8932B2CCF332B2CCCE74359E6984A5B0D2D12B62A652C98D63596323";
    attribute INIT_0F of inst : label is "182490603B332D8D0279838C1CC74143184A58AB9A28842108F2627417608485";
    attribute INIT_10 of inst : label is "32D1D82D58AA4A4D213098572B958843602CE639CC722626692494B203495C0D";
    attribute INIT_11 of inst : label is "495DDC6100AA6D11280D825357ED4BB5CDD2F0E90B481A423A229D699FD56836";
    attribute INIT_12 of inst : label is "B717B03DD555EB9AC495751BCA796012599056CAA1555602DADA23C24AC8460F";
    attribute INIT_13 of inst : label is "AFDD1F597B351240D3484D201E08523105E54FA952B167353393BD719109289E";
    attribute INIT_14 of inst : label is "82DDB36D8C6CF3603BC22AA2A8C22A97F3194631672DB3FC961F2364EDD50909";
    attribute INIT_15 of inst : label is "F6B7DAAFFDFE2AD7EF2E27D55B55EBABE0003FE03FF000FF238D9E008410046C";
    attribute INIT_16 of inst : label is "AABAFBBAFFD4BEEFBBEFD6FAFFFFFE757FFEEB5FFFD4FF53FDFF57FDFEDF77DD";
    attribute INIT_17 of inst : label is "53A55E4900035FFFD9F0038223F3E40183F09FDFA7FE0FFF87B112AAAAAAAAAA";
    attribute INIT_18 of inst : label is "B0000758A240D5649502CAE3122180C3890880B69356894849C96EC063086996";
    attribute INIT_19 of inst : label is "000200000020000000002220431710D9A9B0536C1D19B06D24E24084CA8A6DC5";
    attribute INIT_1A of inst : label is "88888886222108080C401010A4246414840408000000003C16A2A000E0000800";
    attribute INIT_1B of inst : label is "A8A0023400000020424193939090220C86214812521200908111104404C48400";
    attribute INIT_1C of inst : label is "1A0BE736D74FB76C206CCD4AA39CE6F5F9FCFFFF151C451FFC1FF15FEAAAAFA8";
    attribute INIT_1D of inst : label is "C4ED12339A2491058914ADEE7BE9DC93E644E4544D12A64F3D9EDC9940889F24";
    attribute INIT_1E of inst : label is "B034ED29704496EA65AD9ED530097A8AD518A78A14C8021FF7F809A4C9DDA379";
    attribute INIT_1F of inst : label is "273C90D9E34468D20A0F964C036D90069DA2D374DB25B42927B4D399E3EDBD55";
    attribute INIT_20 of inst : label is "874948800160AEDA48D6C167A000E41720025941940A0A2283CCC42CA06A8B68";
    attribute INIT_21 of inst : label is "7B6C52043564A810D4430880D48352412A999616DA883B185283CED50850A92A";
    attribute INIT_22 of inst : label is "901B41069E96C76AB41A9968EC95AC552504854AB2862411004EC0C2941B2B56";
    attribute INIT_23 of inst : label is "337755555555555708421534824729412838E007A44BD710D9018EC302CD0166";
    attribute INIT_24 of inst : label is "38111004F004240000000000000003FFFFFFFFFFF30073007DB4DD5578022333";
    attribute INIT_25 of inst : label is "0920C104190C10480A0014501500A58001003460000140802C801042AE25498A";
    attribute INIT_26 of inst : label is "00C0400040C889027428804002844C006008C880018220104030220001010400";
    attribute INIT_27 of inst : label is "A41145214828A884A422040A5020005000000000000000000000000018000211";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "AC66268BA0A04AAAAB601B654BE6B6AF49DBB9E147C8008106B36D9D2D37FF81";
    attribute INIT_01 of inst : label is "45CA86D5605536A0BAAC04DD413DD626D5A8ED900040A0428008025A9BB994A0";
    attribute INIT_02 of inst : label is "DF52A0996C92FFF49BD40E11D66626093485577552E40923A2EA296A8BAA142A";
    attribute INIT_03 of inst : label is "4B9261A502A29525363403A93066C545214CCB4996A5C270733280804094A0C8";
    attribute INIT_04 of inst : label is "6D2CA068682242CA2D34C0E60380E6020A4D56918652804120824ED499F04003";
    attribute INIT_05 of inst : label is "96880EB1411160880AAC512AB54DB900B414676FBC4E30924A0CF80422449C92";
    attribute INIT_06 of inst : label is "4B41234488B24196908168E24A928894CA924997895D484A0212400862698D94";
    attribute INIT_07 of inst : label is "28C100818203050E80409A412F4006958180B01060203E10235048C1CD9B6836";
    attribute INIT_08 of inst : label is "27E851159113ADA2824AC90440208C8D184841F733512980E313292909529304";
    attribute INIT_09 of inst : label is "0ED54541D74B46968A4A5214A1022449B91BC48929A27A412322448260B488B2";
    attribute INIT_0A of inst : label is "7444E80174A8693AD4200A43A74A4220A23C010009204A6E49B7200350156E40";
    attribute INIT_0B of inst : label is "81146E96A24A0106A10405A00890A42908B4022090A9449011294A8894244AA5";
    attribute INIT_0C of inst : label is "EBFF149128CB764613509A5408B7D00228057B15C42244445530900808094020";
    attribute INIT_0D of inst : label is "545358AAADD0AA17A53A51200208488484169A5D1A94654442974AA94D4CB814";
    attribute INIT_0E of inst : label is "A02510439100808CE320808CD0101518A084052082FA43411290120942518252";
    attribute INIT_0F of inst : label is "F2202068BE0B29AC833B93ADB1E628612148246AB80600000064825D14400915";
    attribute INIT_10 of inst : label is "4EA3537055D49209082412040A0100004C04A5210852C847601894EA136DDD9B";
    attribute INIT_11 of inst : label is "829292C0ED700B93BCD859E3DD87466519C28B070C3820C37A62AE554132F828";
    attribute INIT_12 of inst : label is "6A4813B91113A306292E753814A80D70952AA25AA0AFF01C9493BAC499181B01";
    attribute INIT_13 of inst : label is "6ECE3025514624809400892FE1BC11909A448C66405FAB9329097FFB4080040C";
    attribute INIT_14 of inst : label is "6C9122493171874ECA00310113001136101514A45489B31C02A501292D831815";
    attribute INIT_15 of inst : label is "03400DD555540042AA5555500A90BC5400003FFFC00000FFC3E78DAE906DDF24";
    attribute INIT_16 of inst : label is "035D733000046CCB3282BFAD6AAAA04A06A83500000400100002A15554000000";
    attribute INIT_17 of inst : label is "630417ED000B5FFFDDFFEFBFBCFA17FE7C0F60205000037B8001F08020008808";
    attribute INIT_18 of inst : label is "DFF7FAAEC906DFF100080401804040104204403808870204301080FF10079001";
    attribute INIT_19 of inst : label is "100401151040100000141415AB80201C403880700200401008083F0311100E00";
    attribute INIT_1A of inst : label is "0000000000010100040103006060E0402000000000000003E14052F0C1500440";
    attribute INIT_1B of inst : label is "0A20000100000004060082828180000404014010101000100202000000000000";
    attribute INIT_1C of inst : label is "193C02926134924E5420200F7755A8D1EAF5CFF0105D105FFD1FF11F0222A822";
    attribute INIT_1D of inst : label is "FA5497D3496ADE3B4E38F5AD6BA5F4AB8525A57AA297C5223A1AA511FE0CA422";
    attribute INIT_1E of inst : label is "39C78DD0827F5AB545D40D6AB96FFF8F21593F9FFD748207FFE00103070C52B5";
    attribute INIT_1F of inst : label is "E085FA1FD7BB7508FD143AF8A501DD28D0070950010202F046025A91AF8E31EE";
    attribute INIT_20 of inst : label is "67C98EB6DB73EEDC7CF6E177EDA53D39E9A4D74D74D0CC8BB3ED9C4DA0DE2AC3";
    attribute INIT_21 of inst : label is "432C5A74BD80B9D2D678408CF6F35B91D7D51736DFD33B9964E3CAD651D4B130";
    attribute INIT_22 of inst : label is "F1971349AD36B9997C15A751A93B2AEA49A7E6D33EE7BDA66C8ED1CB271B2B5B";
    attribute INIT_23 of inst : label is "AAAA088282828287FFFFEA410407A6194B6989666773363459C9CDB212CDA366";
    attribute INIT_24 of inst : label is "044A07F0000A920000000000000003FFFFFFFFFFF00010001D575808FAAAAAAA";
    attribute INIT_25 of inst : label is "10022008802260A04011020000000A113260021001580028800147A4014A1241";
    attribute INIT_26 of inst : label is "080100DF202266A480040C20010880208324260080284044AA88800044B44880";
    attribute INIT_27 of inst : label is "84730C084061A881852A444A422053100000000000000000000000000000C000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "011082882222AE38E4A2691039321067FBC884C00257FF7EF92A49040128079C";
    attribute INIT_01 of inst : label is "9CA6041B0730A0D38982724D86449D101C81E62DBB366CDBB36EDB25FF814206";
    attribute INIT_02 of inst : label is "3268D2E68208300EE4412265051034C5A8D12CCCC8EC25984E5824ED3961F68B";
    attribute INIT_03 of inst : label is "34412E673138C68CCDC65A3DCB50B1F1B67324A4681C444718490202AD46362E";
    attribute INIT_04 of inst : label is "18842683191160C11C6C81240C8CA40CE1041A324F0CC92DB25BF106446FBE64";
    attribute INIT_05 of inst : label is "4EF42604C888E26C888E300C617B7AB6766D6B6308C24749636A37FEE9904249";
    attribute INIT_06 of inst : label is "EB0D9CFA9F0D254546D1AF751459E607634D8140E620636318C964486B6D99B2";
    attribute INIT_07 of inst : label is "3DDEC08B9509B326C1B659CE07247D445C3F921F17E6C25CE771A44DA4C76192";
    attribute INIT_08 of inst : label is "9A093C66C8D89C30CB6ECD976412A21DC1BC040D3ECDBE1A78001585C5985978";
    attribute INIT_09 of inst : label is "B071F32E42707160E5694AD2BC99B3248C0950F6CE7B01ADA1A91237C8607675";
    attribute INIT_0A of inst : label is "7752EF9136E30D9B1C9C8B19B3634993599BFEFFDDB6AF3235B994190241732D";
    attribute INIT_0B of inst : label is "101072F2B96258B02594B025C67294A5297C8BB3655776DD8CBD22C473132234";
    attribute INIT_0C of inst : label is "601176E30C0B9B0A48D8431620B912D98685F1AC5E3372232C86DB6129624B13";
    attribute INIT_0D of inst : label is "B7620E08B1120B8CBC8B0EADBD336EB6CEDAC36DD0D753334B5162E73C2EB5C2";
    attribute INIT_0E of inst : label is "E477D9338B2212C461B212C462090C88124210B24AFB6766CE40DB67718A9BCB";
    attribute INIT_0F of inst : label is "083B17641AD1858E38D3495E504680DCA4A437208DF2C6318C66D90073386DC7";
    attribute INIT_10 of inst : label is "B2FB68295ACADEC77B1D8EE379BCDEF6337294A5295B3DF6D6D6622069244A09";
    attribute INIT_11 of inst : label is "31F0F00613FDB901292A0FFB039D52050160F49D10C8C744BA08AEC321944B15";
    attribute INIT_12 of inst : label is "20625F7B2AA8A50D6DFFD2F66A6470975995ED95BA55790EDCD93256FCE8E511";
    attribute INIT_13 of inst : label is "E36FB8D17018F8779197E495E81D2C4C0A4E27D2A10100C945850C58EE76136D";
    attribute INIT_14 of inst : label is "32DDB16DCFFF937379B06F84FDB06FFA50C30420440CB1A2F636BB6DBDCD383E";
    attribute INIT_15 of inst : label is "01000450000155097700000A8E82282BFFFFC000000000FFFC0FEA72529E0E93";
    attribute INIT_16 of inst : label is "89450445C8934110441C3F0500000A022001D4208893224C0000000001000000";
    attribute INIT_17 of inst : label is "01081E12AA040D77FAFFFC7D5F05E801801084080801F800078002080A020000";
    attribute INIT_18 of inst : label is "A0080521F931206EFFF7FBFE7FBFBFEFBDFBBFF7F776FDFBCFEF7EC0EFF86FFE";
    attribute INIT_19 of inst : label is "155401551540155400015400037FDFDBBFF77FEFF9FF3FCFE7E7C0FCEEEFEDFF";
    attribute INIT_1A of inst : label is "101000040000010008000200A020A00280000000000000001EBFAD00C1555540";
    attribute INIT_1B of inst : label is "88A0022001000000020081808180001400004050501010000202008080808000";
    attribute INIT_1C of inst : label is "3008BE590880596CDE3797BA293631196CD627F0101C001FFC5FF05F22AA20A0";
    attribute INIT_1D of inst : label is "C1F2561F2CB924D36ED3A614A592B2A79C95B7D384DE9DBEDD6BB237497BFCE3";
    attribute INIT_1E of inst : label is "D80830A6CD1479AA98A64D545890FA8FFD20F50A568801F803FFFFDBB73C8E52";
    attribute INIT_1F of inst : label is "12C614285D45A8F14982D30341B62AD126CA659B2D82DBA29AD924579096D654";
    attribute INIT_20 of inst : label is "986E7BD96585B123430B0E8816D8E6D736D9713113060120CC10C0148348CE44";
    attribute INIT_21 of inst : label is "CC33A59B4223466D0884A707091C24662ADDE6D9DAA8C466810C3109A47F05C4";
    attribute INIT_22 of inst : label is "1AD340370ADED74A258AD97DB414AD656FB1B866C3D82E40973118340864C424";
    attribute INIT_23 of inst : label is "0001F5FD57FD57FF08421FBEFBFF7CC1F9A2891E188F0EE1624A3C0687324999";
    attribute INIT_24 of inst : label is "02A0800A0020480000000000000003FFFFFFFFFFFCFF9CFF99041D5F78000000";
    attribute INIT_25 of inst : label is "06051C9000800012010E0023E83D500080004001CC0202000000080140108010";
    attribute INIT_26 of inst : label is "F022102014011050008000000010210404900001060003080002508130000208";
    attribute INIT_27 of inst : label is "B24B2CA52B6F9337B5F91839C841182000000000000000000000000002010588";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "420100802626A41040E8000011400247FB8010C2024000000128000D08000788";
    attribute INIT_01 of inst : label is "D8A4744A3721A25B1903720CD70089104803C009B3664C9B3664CA05FF11000C";
    attribute INIT_02 of inst : label is "3470524008203006C0C00265342030C58851288888E805B06C51A4E5B1435299";
    attribute INIT_03 of inst : label is "00810C623110830C8C824A9D8B1221E0972220C08008C00200D12626AC44162C";
    attribute INIT_04 of inst : label is "2A140053199930A19C2C80240584240444001E104E1C5B24B659A0040060016F";
    attribute INIT_05 of inst : label is "CE541602CCCCE16480981024232D3292F22D6A271C4207894328300269800800";
    attribute INIT_06 of inst : label is "E91D15AA95156D4586D1AD75165144078380000240144143308164482924B8A2";
    attribute INIT_07 of inst : label is "188AC0829501932640B6D34A06241544E89287CC22A242CDAF30AC4CE44F2390";
    attribute INIT_08 of inst : label is "0008282708C89890592484B32436C03C88B3B40713CC9C321000348CC488C928";
    attribute INIT_09 of inst : label is "9010A10C4251316245294AD698B1A290820820C004720025B08020036830D425";
    attribute INIT_0A of inst : label is "5362A59032410599181C8109932381B75B1800003CB62F22B491143900C12224";
    attribute INIT_0B of inst : label is "901022509322489024B49024C65694AD6BFC89917055364D8D9D224473176234";
    attribute INIT_0C of inst : label is "4022727208091C1A49484912009112490685E8A89E3122236C96492369204917";
    attribute INIT_0D of inst : label is "933204089116098D9C891AA4953B26B24ECA4934B0534333495122673CBAA480";
    attribute INIT_0E of inst : label is "E477C831832636446196364472191C8832C631965A792F22DE404927319E9959";
    attribute INIT_0F of inst : label is "201B57441A4115081153017C70860048A5C4360115E2421084624808336F64C7";
    attribute INIT_10 of inst : label is "B24A0929CACA4EC67B1DCCE371B8DCF62276B5AD6B4A3CF2D2D5006100008809";
    attribute INIT_11 of inst : label is "31F0704003FCB840420007F90911424D03605095008804409A28AEC2208402F5";
    attribute INIT_12 of inst : label is "24405CD92AA9362624FFD3BD2ACC200748B1E0151A55790E4C48444278884700";
    attribute INIT_13 of inst : label is "E378A9D33218FC738196E49F200FA800021A0862A0204480EE6E34096C56026C";
    attribute INIT_14 of inst : label is "224C91248FFF9323F9B00F80FFB02FFD50460420440891A6621399249CC53C3F";
    attribute INIT_15 of inst : label is "AAAAAAAAAAAAFFC082AAAAAA0AA2A88BFFFFFFFFFFFFFF00000B0160EF0F0616";
    attribute INIT_16 of inst : label is "AAAAAAA82088AAAAAA82AAAAAAAAA1B08EA82A28A0888222AAAAAAAAAAAAAAAA";
    attribute INIT_17 of inst : label is "03000E24FFF8F28804000002800810003FE0002053FE03FFF849E2AAAAAAAAAA";
    attribute INIT_18 of inst : label is "00000081000EDFE000000000000080008000003000060000200000C000000001";
    attribute INIT_19 of inst : label is "140154151415415400000155AB00001800300060040080201010000200001C00";
    attribute INIT_1A of inst : label is "10101000040100000403010060E06000020202000000003FE14052FFD4005540";
    attribute INIT_1B of inst : label is "2020000A4040AA080A0282838280401400004050105010000000008080000010";
    attribute INIT_1C of inst : label is "3008BE4B0180CB68CE1793B26A72130BA46267F5451C451FFC1FF41F88020208";
    attribute INIT_1D of inst : label is "91F6549E2CB984D26ED32235AD32A6A535951F13805C98B0503992264163FCE1";
    attribute INIT_1E of inst : label is "681C1682C8547B001C06CD00E800F28FFD20F50A562003E7FFE003DBB7380E52";
    attribute INIT_1F of inst : label is "10C6A4301E01C0010986D10101B2880382CA248B6D825BA69AC9305710926340";
    attribute INIT_20 of inst : label is "00682BCB6F05A001D39E0811125AA2C5164930010004010048E0081808440608";
    attribute INIT_21 of inst : label is "C000041800000060000CA0060018002C2A888271CAA8802000188000243C0504";
    attribute INIT_22 of inst : label is "1AD1023582DE4542017A59250415E56527B19E267BCF2E429720180000C00000";
    attribute INIT_23 of inst : label is "AAAA2A088A22208FFFFFE08000077C80F892801E10070EB100001C0684004800";
    attribute INIT_24 of inst : label is "691407E07010240000000000000003FFFFFFFFFFFFFFFFFFF90410207AAAAAAA";
    attribute INIT_25 of inst : label is "881842056549104C0CC04418044000840198A5001080C8062410201006206082";
    attribute INIT_26 of inst : label is "0400201F4100810B4B20B01004C5001A004801560182A88050200800020A0000";
    attribute INIT_27 of inst : label is "924269AD6B4F11171CB91C7BC861083000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
