-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "29127CAFDF5829A327973996FBBBBB09EBDECBBECA5A0A56B0FA063608A4922E";
    attribute INIT_01 of inst : label is "F1DC3D67BD91CE3B87D891EE4F77207DE341A5C6F0D2EDE5B96C3B8DB7FBD29F";
    attribute INIT_02 of inst : label is "9DCFDEEFE772DA3489E4299CDC43CEC3B0DBDBB0B623C6D347F0CFFB696DBBFD";
    attribute INIT_03 of inst : label is "66412F9CBC191BFBEFBEFB26364F78364F604BD8F6E4EC6B96CF9996E73F7BBF";
    attribute INIT_04 of inst : label is "36F6E3EF98C004F5BDDE0C1C7690FC60633217C6430DFE6FF204E6C7E119FB98";
    attribute INIT_05 of inst : label is "10F8780299949C91979F7DE5B2DFAB3CF7B8E99823BFFDBE2DFC9B8236764022";
    attribute INIT_06 of inst : label is "2D9707693E3FBFDADAC0323B1F9B9BDB9FDBC7E100123A4CC4CC077BDBC00002";
    attribute INIT_07 of inst : label is "B726B3642B74D66C8EB7C99B026D34997BF0110C800939391FC01DB764E7B977";
    attribute INIT_08 of inst : label is "6D1D0AAE4B95BC992C844CFB8D6D1956D15BF10FDB9359B26CD675BA66C8C424";
    attribute INIT_09 of inst : label is "7FF7712ADE03E35A7FBF5BC5B5E25CF9835D5541406AAC1B45A8E82616ED974F";
    attribute INIT_0A of inst : label is "F4B7FEA5417FE5D97FEE5CBFF72FF765FEA5BA97FAB7FF7FF777F7FFFF777FF7";
    attribute INIT_0B of inst : label is "FAA5AB427FD4A96FFDCBBFFF72EFFFDF4B24D25B3FFFFEE5FCB7FEE5FDB7FEA5";
    attribute INIT_0C of inst : label is "EFFEFBFFBFFFFFBEFE0072EBBFF72CDBFF52AFFFD4ABFDF97F2DFFB92FFDDB97";
    attribute INIT_0D of inst : label is "BFFF6DBFFBFFBFFFFFFFFFEFBEFFEFBEFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFF7FF7FF7DFFFFFFFFFFFFFFFFFDF7DF7DF7DF7FFFFF7FF7DFFDFFFBFFFFF";
    attribute INIT_0F of inst : label is "FFBEFFEFBEFFEFBFFBEFFEFBFDFFFFFFFFFFFFFFFFFFFFDFEFBEFBEFBEFF7FB7";
    attribute INIT_10 of inst : label is "05042020420A52804200058F2F3C3E3F1FD8FA16F8ADFFFDFFFF7FFFDF7FF7DB";
    attribute INIT_11 of inst : label is "E48DAD6A5296885179F9E20CE7EC0F803E01F00F8003E01F040F80101F88404A";
    attribute INIT_12 of inst : label is "3F800050C3CDF997B5CE8EA345EF29997A631F8FC3E3B1F8EEDE80C062104263";
    attribute INIT_13 of inst : label is "4204247DD93E7A267EF439DEBD79B8EED004044106010042000FFC0040000882";
    attribute INIT_14 of inst : label is "F7B8DC63E1FF60DE68C4082123F0FD8FD9FA3F1FDA1266141E5222F914A5294A";
    attribute INIT_15 of inst : label is "8D13098EC7E41B36DCFCF7A6F48FEFEDBEDB98F304C51A47E1B1F8FEC5B6E424";
    attribute INIT_16 of inst : label is "731E61314691F87C7E3E2DBD9E00C1884482208250A0810408414A50084020A1";
    attribute INIT_17 of inst : label is "14D45D3738FC761F0D8EED09044101285040820420A528042010509C7DF6DBDB";
    attribute INIT_18 of inst : label is "0C030040303E000000000001181FF8104004700401E0102F84C39B113F8C30C3";
    attribute INIT_19 of inst : label is "12492DDB3A686E6F33A9F774C89DCEFAE338EE78C9A45FD63528984D99FCE000";
    attribute INIT_1A of inst : label is "C43F377BCBD7E2DDE9B313C49D00E60180005C7F594DB3739E0A3FC688EED873";
    attribute INIT_1B of inst : label is "6EF96004DB3D0F9B264F82443B5300011000109A7379F4347F3B8C9BFC43729B";
    attribute INIT_1C of inst : label is "DA7B9B1FFFFEEADEAD0AEF7BDE46F6779583F8842B68B5F4BCCD65E7375A7A93";
    attribute INIT_1D of inst : label is "77A37BDED4DD3B27492792F59DC77E777587EFEFEF6F6A5B3CC3CE1D9999CD39";
    attribute INIT_1E of inst : label is "3C6D4A138AC7F9AF9C724DD21DC349490E18394F4E48FEE7B52BA4B3B7348CCF";
    attribute INIT_1F of inst : label is "1BCDDDDE97A0DCB5CC9E632B2BC2F74A256DCD3BCCEFF5D1DA98D4C6E1CFCC7D";
    attribute INIT_20 of inst : label is "6C783FE76B1C925D3DD89CE5FB5BC78EC7E6FDD1C3C44A27FFE63F429E833E33";
    attribute INIT_21 of inst : label is "32FB5BFFAD5E750F7ED1FF517C07B7F3CF5DF27BCFCAFBBCD49A76D23478AEAF";
    attribute INIT_22 of inst : label is "DFBF7EFDCFBF7EFDFBBAFEEFBC542CE73DCE604FE627A7D01DE5E545DA848B77";
    attribute INIT_23 of inst : label is "F7EFDFBF73EFDFBF7EFDFBF6FFFEE003F9FFFFF7F3FFF3FFFFEFEFEFEFE7F359";
    attribute INIT_24 of inst : label is "FEFCFEFC7EFC76EDDBB76EC7CF9F3E7CF9DFDFCFDFBF7E3FBFBFBFBF9FCEFDFB";
    attribute INIT_25 of inst : label is "F1A9FFFFFFE7E7F7E7F7E3F7E3B76EDDBB1F3E7CF9F2FFEA8FDFBF3F7EFDF8FC";
    attribute INIT_26 of inst : label is "DFB5FFFC7FFFFCFE6B7FFFFFF9FDFDFDFDFCFFFCEFDFBF7EE7DFBF7EFDEFABF3";
    attribute INIT_27 of inst : label is "8E5D7BF6F76DCE6E3DA03F7EFC7F35BF7EFDF8FEFEFEFEFE7FFE77EDDFB9F7E7";
    attribute INIT_28 of inst : label is "69B50DD37300FB979E38C8921DF3E6461710A8B264C9938615FDBBD7C772DE5B";
    attribute INIT_29 of inst : label is "D6687FCE13873A43691B18E50C7FDB8142A6E9AC03EE5A18999A84F305390129";
    attribute INIT_2A of inst : label is "B7EFBEDDE3BDEBEF1A70EEEFB7D657D7AF965E5C7F7FF6BFA668F3272069E786";
    attribute INIT_2B of inst : label is "53F8FF8EC7D8BF667D8BFE71FC79E1E3FE2D999FCBBFBFC0861F3B9BE336F9CD";
    attribute INIT_2C of inst : label is "5A0977FFD1111112C65669863B4E1DC49D385F3A447E3F1FFFFFFFFFC4444D3E";
    attribute INIT_2D of inst : label is "F1404A00FBCBF22CB80F4FA4A7252BE237ED9633FEA00A58C8D9381099161F41";
    attribute INIT_2E of inst : label is "1EEDBCEDD7397A5CDDDBDEB7ADC77B9EF0EE8016A104FE4443CF120AA997A722";
    attribute INIT_2F of inst : label is "9C773EF997D38FCF1EDDE7F4DB3F7BE2FDB1A7D9B2367E7B0F73ED5A919F47A7";
    attribute INIT_30 of inst : label is "007E1D77DDF77DDF731AD6FBEB17B13CED34E57B3FD3958DD6FDC779797C597E";
    attribute INIT_31 of inst : label is "00050664000000802FC800000AAAFC00181100A09000000080020F00001F8000";
    attribute INIT_32 of inst : label is "04016900011504447840001800282B1200030000541190000020200000800000";
    attribute INIT_33 of inst : label is "01660000000156BF8000040802228C000050005057E00000000002B820002804";
    attribute INIT_34 of inst : label is "0055F90000002A29E200058282A120007E00000501000180000A2FC800011100";
    attribute INIT_35 of inst : label is "BFFAAFF000F0008007C8001F800445244000FC002220A2000002AA8020000800";
    attribute INIT_36 of inst : label is "FF5D7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA";
    attribute INIT_37 of inst : label is "7AF3D924FCF0023D98F7ED3CE9EDEDDE7B2DB9E04040937A8DC6C8A7F83FFFFF";
    attribute INIT_38 of inst : label is "31BF9EF9E4EF79329CC8E9A8B73F9E44E3F57B7E7C3E1F1FD37F9C75ED4DFBBB";
    attribute INIT_39 of inst : label is "DF3D3AD8925C8DBFADC43379E7CC83DF3CFDECB9BE7DEF21FCDB5E79FBDB8FCC";
    attribute INIT_3A of inst : label is "4402094282020420A5280421510423C001040FECFBB3EECFBA5AC27CBDFCEB7B";
    attribute INIT_3B of inst : label is "8D9CFB93699642A0733BBBF8E1782FD805ADEF98F7CEE1EF0B179F8CF8EED004";
    attribute INIT_3C of inst : label is "010200000080000000075F846B2C04D702162C59DBF66B7B0E7CDF39B791BB9E";
    attribute INIT_3D of inst : label is "0045000800000001544000000000000000000000007570000000020000400080";
    attribute INIT_3E of inst : label is "02100210011040088800882108C6398E7403F90826374E561004000200000000";
    attribute INIT_3F of inst : label is "E10F7D74A6FCE10F7D74A6FCDFF7E87FE400700E0380701C1108011010048100";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "000080102CECEA5CD94F6F4BA84446D63E232CCB2AE8AFB0CF6BD512A69DD802";
    attribute INIT_01 of inst : label is "0B5505C4EF4F1FEEA1700830209D28C396F29A3DD94C1BBA7C380883492C0C60";
    attribute INIT_02 of inst : label is "4325018280C02C9923B11C0A2AF1233841022ACE6977D82529181492DCDA4882";
    attribute INIT_03 of inst : label is "551852214628804EB90954CA18018C18018C056819B03A2483013A895004864A";
    attribute INIT_04 of inst : label is "8D1928D78442C07B4331835D61A313D969EECC20B48AC55628E21B189CA118E6";
    attribute INIT_05 of inst : label is "1D4EA67E24F22B222A69E64A65A0541179E64C6029461A49922675F8C8AC8FE0";
    attribute INIT_06 of inst : label is "1259ECCE59E6E873B38FF3A9D4F8FA30FA264FFFFFF3A8A8A8A800A6747CFCFE";
    attribute INIT_07 of inst : label is "4BCD6DD406B9ADBA844B336E81201498AE755ACFC40AEAEAE27C044F89634088";
    attribute INIT_08 of inst : label is "B7C865D1A5AA5E100880261250974C897AB5F50DA5E6B6EA05AD4A5CDBA820DB";
    attribute INIT_09 of inst : label is "088000012F004CB24644A5FA42F803877EA80280155D595FE6555799245381D0";
    attribute INIT_0A of inst : label is "F6FFFEB765FFE774FFEB76FFF5BFF5F3FEF3BBDFBB7FF88988B9810228000010";
    attribute INIT_0B of inst : label is "FEB7E7DB7FD6EDFFFD6EF7DF5BBDFFDFEFB7FB7FFFFFFEF7FE6FFEF7FF6FFEB7";
    attribute INIT_0C of inst : label is "2000000001001000042D5BBDF7F5BBBFFF7BFDF7DEFF7FFDFF9FFFBFBFFDFFDF";
    attribute INIT_0D of inst : label is "4001124104104100000124000100000100000004000000024900104100000000";
    attribute INIT_0E of inst : label is "0000000042080001002018282002080002000043043000001242000000410410";
    attribute INIT_0F of inst : label is "000000014414510514414510530820861861C618608208082082082082048068";
    attribute INIT_10 of inst : label is "FDE7FFFFF2FBDEFFFE3FFC3301CD0A8150AFA9C19EDBFE800820020000000000";
    attribute INIT_11 of inst : label is "1A33BDCE7D2A440DEC64D5605924FF9FFE7FF3FF9FFFE7FF3FFF9FFFFF8FFFFB";
    attribute INIT_12 of inst : label is "3F8FFFC821FF1FC1843FC15458171C0A009150A150385D0A953BE7DFEFF0A03A";
    attribute INIT_13 of inst : label is "5FFC0F428170B692E36DE0754A970A857CFFFC7FFE39CFFFFCFFFFCFFFF3FFFE";
    attribute INIT_14 of inst : label is "DA7BA7746DA62C6678E5FFE07A1426A36A06E156AFAEA037EA5FE2FF1CE739CE";
    attribute INIT_15 of inst : label is "0BC880E3742DF69DB7631FF18B7276D653AC542A403454742A946AB57EC93A09";
    attribute INIT_16 of inst : label is "8A85500D151D0AA51AADD24AF7E7DFBFC7FE3FFFDFBCFFFFFE5F7BDFFFC7FF91";
    attribute INIT_17 of inst : label is "3E3E02431E85028542A957CFFC7FFFEFDE7FFFFF2FBDEFFFE3FFC8E187CD4635";
    attribute INIT_18 of inst : label is "FC3F0FC3F0FE3F0F0F0F87871FFFFFF07FFFF3FFFFE3FFE047A0E1C011000000";
    attribute INIT_19 of inst : label is "4D36D274EAEC999A6C5408FE13223BA3BCC619D456D542A3AEFFF080FC4FF3F0";
    attribute INIT_1A of inst : label is "BB4CC286E6741983FC6DED3A473FFE7F9F0FC789E01F66C2624281216A95771E";
    attribute INIT_1B of inst : label is "D5041F5A4613846C09F0086944AC3F3FF1F9FF84E514D54A8CCC22388B541F3C";
    attribute INIT_1C of inst : label is "719C76E24A491F29F04118C631B1890C48CC0718D6C142F80232D2585470A54D";
    attribute INIT_1D of inst : label is "DC70CCB1FE378D05A58F6C9E3632CC8D9F50FCFC17B7B50E9082AB871514DBE6";
    attribute INIT_1E of inst : label is "E297E9A8602206013E5D3DE3121CB6A5A34D4CE63B29930F7A965AA8E8C7CA82";
    attribute INIT_1F of inst : label is "FD663221447F12E4B269B600D5B50BB4A0C6A2AEA0326E3E75544A2A3BAB20D7";
    attribute INIT_20 of inst : label is "FA975C5966E33537CA372D6AE4ABA9793C7865BF7C13B4E890C9F33B43F491F4";
    attribute INIT_21 of inst : label is "CB5625BF8AEBBE18017A7BEEFE004C87B04755A4F120256F2B4FDD7C92941119";
    attribute INIT_22 of inst : label is "24509102706281820615512FD78C5296A3AD313050DAFC7F3332513A263B0049";
    attribute INIT_23 of inst : label is "091024409C103040C103040EC0C100240B0200181400040010383830382914AE";
    attribute INIT_24 of inst : label is "0103010281018812244881182060C1820541C1D000000040C040C040A0310244";
    attribute INIT_25 of inst : label is "8A56000000080808080804001C48816204E0C10B040FC0EB9010004081020503";
    attribute INIT_26 of inst : label is "B154157681820520948000000206020602050203102450911820628182A0AAE4";
    attribute INIT_27 of inst : label is "66B49CDD99961DBEA4CF408102904A40000001030103010281008B142C522C50";
    attribute INIT_28 of inst : label is "F1D9CFE9BDFB5DE604022025F7C98DFBE047B5B13B74ED73EAE2EE3C3CCDB1B6";
    attribute INIT_29 of inst : label is "2A96811EFDF9CA2AFED7E73BF7DBE4FBA7456497ED779C674CACE5EDF38E6ECC";
    attribute INIT_2A of inst : label is "D9BAEB82008385E2E59311104D3DABEE786D35B312592D4970882898D15E9849";
    attribute INIT_2B of inst : label is "1DC449400B352CD43340C51D3F0CF8F8C202EC47389C8D40ABA3CEE4D9FF477F";
    attribute INIT_2C of inst : label is "B0969E1E1555555411195B15CEB382C86EDF31DFB74FA7D3C6F3800B00012BDD";
    attribute INIT_2D of inst : label is "A55031E117A7EDD7DFD0E25A58C0801D9C9B4D8D18AAAA0222BEEE464CA76012";
    attribute INIT_2E of inst : label is "67BB6F3B3C79D221E7768EE3B37233744A1B3C25C9C15FFB3C30CCBAA089C1D7";
    attribute INIT_2F of inst : label is "3FD96B874D27F1F6CBB6593C24C79ED92740DBA610EDEFC4A1C5B9F1CC2DF2FC";
    attribute INIT_30 of inst : label is "FF81B77DF222A08288F39C5924E844C1985A3280D528EA436D76ED058ED3B4C9";
    attribute INIT_31 of inst : label is "00787E7DB001010000370000040103F6E6001806002FD40000C0000B64BF8007";
    attribute INIT_32 of inst : label is "002002AE2000200981997178010140CDF8098001028072D940000333FF965A00";
    attribute INIT_33 of inst : label is "FC19E3E0E0010000001BD0200DEC20B64AA00068199AB8D08002BDFCFF909440";
    attribute INIT_34 of inst : label is "1AA1C6E400A940004E4000034A8CECB682131001F76E3470004900342DE80010";
    attribute INIT_35 of inst : label is "BFEABFED84F0A08000F725BF80000029E96DF802400955400003FFC0C4978800";
    attribute INIT_36 of inst : label is "880340AA97D40FF83FF96FF297F32BE455D9AA37C00FE83BF1655280030004EA";
    attribute INIT_37 of inst : label is "CB082CDB33104382E3193877A75B5A6105D2674040C19B7EDFCB718DB3D10025";
    attribute INIT_38 of inst : label is "0F6EF3275389C4DC7327A757CC7371339CD9CCD98D0A8142255165435712084C";
    attribute INIT_39 of inst : label is "3CC205BC6D203264FA602C8810387644CB3A3440C9C1389F77AE6196644C1B2A";
    attribute INIT_3A of inst : label is "C7FFFF7EF3FFFF2FBDEFFFE3F17FE3FF3FFC11B14EC53F14FDA739504A0016E0";
    attribute INIT_3B of inst : label is "BB4745B6B6E817C0CDCECE8C1CCC8417801A334338A5CA71C68804E20A9573FF";
    attribute INIT_3C of inst : label is "AD5AAAAAAAAAAAAAAAAD770195021C3D0E2902A244D934BEED8FE8EFD9B654E6";
    attribute INIT_3D of inst : label is "D555556AAAAAAAAD5556AAAAAAAAAAAAAAAAAAAAAADDDD5555555AAAAB5556AA";
    attribute INIT_3E of inst : label is "FFFCFFFF3FFFF3FFFFCFFFF52DEA5A9EF4FFFFFFE54FE2E5555555AAAAAAAAAA";
    attribute INIT_3F of inst : label is "2153CB8B5D12E153CB8B5D12E5389F8B3B9FF3FE7F9FF3FCFFFF9FFFFCFFFFE7";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "A83EB6BED910C0208FDAA11D1C0003E800024B65BAA09D244F8193D9FA9934D8";
    attribute INIT_01 of inst : label is "8E626BF960B2D1EC4DA7D6DB5AEC4FD6263FE5190EF3821F21D2EE7A5B4F77ED";
    attribute INIT_02 of inst : label is "97CFEBF5E5F32CD9723EC375950CD598CFA7D566798828740CE3792017924C01";
    attribute INIT_03 of inst : label is "FF9E58216BF636B659FE3FC9E99A97ED9ADFF7B9A98F537CED1A75ECFDEFAFDF";
    attribute INIT_04 of inst : label is "D9A929F8FF2D5B42C626746B47AD3F65D8CEBFFF5F7A18D0C4FDA529F7326333";
    attribute INIT_05 of inst : label is "FD9EDE6F2BFFB7BD47D20987D37FAFE53B7A5227E88002D69FFCB27DCEDACF2C";
    attribute INIT_06 of inst : label is "FF2EFCD14C2BDFF5864A77DFE9B5B5F5B1EC8FB91387F37777FFF41BA4BC30CE";
    attribute INIT_07 of inst : label is "F4D73C78DF4AE78F19F4F5E3FF6D3043408828137DF737373FBFF762F352FFFF";
    attribute INIT_08 of inst : label is "D9E1F00E7A47A36051117727E3EAE23EAC7A0A3A7A6B9E3C18E7F7A578F1FBE1";
    attribute INIT_09 of inst : label is "CCE44457D1FEB80DBB9B7A3075096D9B7FD7777E9A8806AB58082FC4C8BC463F";
    attribute INIT_0A of inst : label is "C0D379762DF7963DEE9762FB4BB54B347D65A4DDA47DE4CBCC776D46E6CCCCFF";
    attribute INIT_0B of inst : label is "5B37CFBFCEE6DDFFF248A418B2694E3CEFFE9BDFAE1F7937C4F77D37C5F73D37";
    attribute INIT_0C of inst : label is "B65B6DB6DA6D965A6985FBF3F8FFB9FDBCF2FBCF34AA533DF734CF7FBCBF1ADE";
    attribute INIT_0D of inst : label is "9B6D925965965964965925A6DA6DA6DA6DB6DB69B6DB6DB6DB6DB6DB6DB6DB6D";
    attribute INIT_0E of inst : label is "4D34D34D75DB0DB3EB85BEFB4D34DB6F3EFBCFFFFFFFBCD37D3EF3EDB69B6DB6";
    attribute INIT_0F of inst : label is "BEFAEFBFFFFBFFFEF7DF3DF7CFF38E3CF38E78F3CE38F3EDDF7DF7DF7DF0879F";
    attribute INIT_10 of inst : label is "29E2FAF7501A1E9A640C3D3DCA35769F4F2F90CDA7DF797FFFDFFFD77D75DF5B";
    attribute INIT_11 of inst : label is "3EAC044B5422A9AE83BAA27B6654FF03B429A1BF1243C27A35ED03DA5E05FBD3";
    attribute INIT_12 of inst : label is "1983A85BCC50EA321E42A80AD948636AD6ED59A5D6FB3E9A59236794CBE74DBD";
    attribute INIT_13 of inst : label is "1AF5EFA7A77B2EEEF45DFB3F7EFFFA596CEF587BDC010A775CBFFECDFD33CB88";
    attribute INIT_14 of inst : label is "184F23FC2FFDAFF050A06CEF7D3669AF9FFF9F4F2DF37580FC1320F814E7394A";
    attribute INIT_15 of inst : label is "365136FDFA79E69D120DE4ACF7314B25264F89B11B3A7DFA6B74BA4978DB9EE9";
    attribute INIT_16 of inst : label is "F13626CE9F7E9ADD2E9796E2F1E78F2F80EC1BFA9E3C2DDEEA0343D34C81BBB7";
    attribute INIT_17 of inst : label is "018190BE8F4DFEBB4FA796C1A029EF4F1E16D37501A1E9A640DA5B6D60727089";
    attribute INIT_18 of inst : label is "EC070D42F0FE140E010D05870BFFFBF03DDEF0772FC0D3AEDB4DFFBE8CE49249";
    attribute INIT_19 of inst : label is "E9B4D3665214CED147036815B3BF7B810B46BE4F13755FFFCBC27F7DA39B1250";
    attribute INIT_1A of inst : label is "10C66CED6A6C69612B117AD7C61FA63F96029F8266D249590D36B6CCDA59632D";
    attribute INIT_1B of inst : label is "58DB3402BAE3AF94FD1FD719EE841F3DC0F89EACD6D42D27976E7736E0D25DB4";
    attribute INIT_1C of inst : label is "92DFB06C4C46023023E1000000CC023092D026420382251343F026854C97C09A";
    attribute INIT_1D of inst : label is "E557076681C0719A5EA95721D9C1533221831B3818998252E6694459D9D9386E";
    attribute INIT_1E of inst : label is "0C4822D620379442B2E2F12D7C782B4E8104212BC158AE6941616711254B5CED";
    attribute INIT_1F of inst : label is "33DC88DA9784316F742C24848A38945DF319CD72CE6ED1C396B995C49E46CE48";
    attribute INIT_20 of inst : label is "0B91A7A2583C4AF83DC15AD59A52C6969D89B8438E25CA8DAD36468CBC0B666B";
    attribute INIT_21 of inst : label is "D1BBCA006405C4977EB5844701F5B574A0A92A598697FBBB04FA2487646F406E";
    attribute INIT_22 of inst : label is "F7FFDFBF6EDFBB76EC955056C06384E72D4E5E5FAFA50183D5782E5801ECEF32";
    attribute INIT_23 of inst : label is "F5EBD7AF53A74E9D3A74E9D3959523EBFCF9FFFFF9F3FBFFFFF7FFF7F7F7FBDD";
    attribute INIT_24 of inst : label is "FFFDFFFF7FFF7DFBD7EFDEB76EDD3B76E96B6BEFFFFFFFBFFFFF7FFFDFCEBD7A";
    attribute INIT_25 of inst : label is "FDEDFFFFFFF7FFFFEFFFFBFFFBEFDFFF7EDDBB7EEDDBD5EA87FFDFBFFFFFFEFF";
    attribute INIT_26 of inst : label is "EFC2AA823FFEFEFF7B7FFFFFFDFFFFFBFFFEFFFEFBF7FFDFB76EDFBB7605055B";
    attribute INIT_27 of inst : label is "A4F1946909C090B2892F1FBF7F7FBDBFFFFFFEFFFFFDFFFF7FFE7FFFFFF9FBF7";
    attribute INIT_28 of inst : label is "0F685B797C728248DFA62730EA5948B8CF01D4418A16247085354C4DC88BFFFF";
    attribute INIT_29 of inst : label is "35068021E23044C1DD0EDE086B30003BE7BFBCF1CA0927EB4CB42DBC70D4E9D4";
    attribute INIT_2A of inst : label is "485A95101C215A2DC0C0800006C814F09989FB7D201240120DEEF898DE3E1049";
    attribute INIT_2B of inst : label is "FCBFBEFAF04A09A186B29A549563BF3B3DBBA5B8343EE94FAFE456EC29ED127F";
    attribute INIT_2C of inst : label is "00D6EE667FFD555F31323FE3D415D0BFBB77DEE33FA399C8EDF3FFF87F5607CA";
    attribute INIT_2D of inst : label is "EF5FFBFEE95950CB21EF67A5A19B77A8C9E9B4D92BFEABE6247C77CA6EFDEF12";
    attribute INIT_2E of inst : label is "C1A921511564498126221204840040809A7CBFBE7AFEA191397F4FFAADED7641";
    attribute INIT_2F of inst : label is "B398C5DBC47672A94DA658E83FCAB7290B77FD407DA5D10A06D6E00210A60100";
    attribute INIT_30 of inst : label is "FFFFD7F7D20A28755C9765555B97997EAB45B06EE213C1BB9281B84237EDFC53";
    attribute INIT_31 of inst : label is "FBD7D7E44C0FFFBFE85AFFFFFBFEFFC97FFFEBEB9F3B5BFFFBEFFFCCD3407FFF";
    attribute INIT_32 of inst : label is "EAFF7D2B7FFFF9DBFE457087FFFAFE1FB8171EFEFDDF91B4BFFDFBBBFDEE459F";
    attribute INIT_33 of inst : label is "2BFFE697FD55FFFC711AAFFEFE1CBCCE4157FFD7F43DCDEFF75FEA3DAB917FFE";
    attribute INIT_34 of inst : label is "F5551FD1FFFFFEABD2AFFFF8B56773487FFFFFFF0112380DF7FEA218AD5FFFFF";
    attribute INIT_35 of inst : label is "141414110BFF7F7D5FD8DA407FBFFF8345DA07FFBFFE1AAFFFFC003F2FFD47BE";
    attribute INIT_36 of inst : label is "FFA57FFFE3D6A2F97FFB7AF43D763EA75F57AF03C363E871F170583AB67FEF14";
    attribute INIT_37 of inst : label is "D58A05F73907C4A0770FD6679B16B3B140F6DA479F1DDDF1BB7C87224BDF8FB1";
    attribute INIT_38 of inst : label is "CE6F374D634248FBB747320AD946A23DBCBA97D5952E934B749CA52F16DE0207";
    attribute INIT_39 of inst : label is "0762A1675FE732613B37EE954290FEBAC5264B49D358491B79BDA58A4C949ACC";
    attribute INIT_3A of inst : label is "C1F6DA78F07F7501A1E9A641415FE3DF21E1FACE944A552955F1FF47F6028582";
    attribute INIT_3B of inst : label is "334A666CB36D124486D4E6718CD62E4FF7FA10B70D5D0E5AF9785A6EBA5960DC";
    attribute INIT_3C of inst : label is "F7EDDDDDFF577FF9FF7D7F7BC7D0401E2041D319DBADCF42F397B74F687FBF30";
    attribute INIT_3D of inst : label is "FCBAF2FF7FFFDFDFFEFBF7FFFDFF45FD883E79E79DB5573FF5FFEF9FFDF33FDF";
    attribute INIT_3E of inst : label is "DFD43BDB37F7504FFCC2FF9090A429400057FF2A0DA15AB3F3E7FFFE7FC5FDFF";
    attribute INIT_3F of inst : label is "9F72C4810D049F72C4810D04AB4B28FAE7888310481000C03F4893B3D435CBA0";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "AB937EAFCF7CABEF77B7F7DD5BFFFF8BE3FEEF5D4E56447670FA33AFF9B23ABC";
    attribute INIT_01 of inst : label is "7BF97DEFFF87EE7F2FB8D7D75E6BA0E8F741A5F2F0D2F5E5F5547F09A7FF52DF";
    attribute INIT_02 of inst : label is "DDEFFEFFF77ADA348DC6FB89EDDFDD6FD17FDF5BBA67C49B6AFBCFFFFFFEDF3F";
    attribute INIT_03 of inst : label is "6EE13D9CFC15BFF7DFBDFD362F5FF82F5FF06BD1FFD4DC6FD5DFD9D77FFFFBFF";
    attribute INIT_04 of inst : label is "5FFFF5E6CEB7BFF0F7FE0C1677D3FCE0337717C6A38CFEE7F704E55FE97DF77C";
    attribute INIT_05 of inst : label is "1AFD799099D7DFD1BFBFFDB6BB5AFFBEE73BE4E833BDF6DEF6EEBF827B7B7892";
    attribute INIT_06 of inst : label is "FDFE0BABBEDFDFE9FBF14B7BBDDFDFEFDFFD73CA350B7EC44C4407FDEFC3FF0D";
    attribute INIT_07 of inst : label is "FF2CE3467DF59C68CFFFCB1A0249B491EEF2FBA0D40D7D7D6FC03FBBBFFF3FE7";
    attribute INIT_08 of inst : label is "67793F7EEFFEFF93A8CE7FFFBDFDFBDFD3EFF38E7F9671A3699C6FFAC68CCEFE";
    attribute INIT_09 of inst : label is "F77FFBBF7E07E7F83F7EEFCFB7FEDDFB83FFFFC3EEEAAFBB43FB78267CF7BFDF";
    attribute INIT_0A of inst : label is "0902105A92008A820081A10042D400080049402041800777777FF7F777FF7FFF";
    attribute INIT_0B of inst : label is "045A02108403468D20344BA02D52E000B449AD806000005B0D02105B0C02105B";
    attribute INIT_0C of inst : label is "FFFEFBFFBEFBEFFFFA5C0D12E900D200040D12A00344B816C34084145408006A";
    attribute INIT_0D of inst : label is "FFFFFDBFFBFFBFFFFFBFFFEFBFFFEFBFFFFFFFFFFFFFFFFDB6FBEFBEFFFFFFFF";
    attribute INIT_0E of inst : label is "FFFFFFDFFDF7DFFDF7FBFFBFFFFFFFFF7FFFFF7FFFFFFFFFDFFFF7DFFFFEFBEF";
    attribute INIT_0F of inst : label is "EFFFFBFFFEFBFFBEFFEFBFFBEFFFFFFFFFFFFFFFFFFFFFDFEFBEFBEFBEFBFFFF";
    attribute INIT_10 of inst : label is "429B45109D452D0E11E6033FAFBEBF5BADD1DB7F78E001FFFFFFFFFFFFFFFFFF";
    attribute INIT_11 of inst : label is "E68D296A5AD6ADDB75FBF37EF7DFA2F38BCA5E42E0A0BCC5C8B2F1A9C5769915";
    attribute INIT_12 of inst : label is "FF7160386FEFBD9FFEDEB6AB67FFFADDFF4FAFD7EFF5BBFD6EDC192298A86BF7";
    attribute INIT_13 of inst : label is "A45A26FDD9BE7B2F7EF63FEEFDFAFD6E83023B8009C632813B400332340E2541";
    attribute INIT_14 of inst : label is "F7B97867F3F770D9B77A019137F16D96D9FA3FADD01266A31DA11D00EF3BCE73";
    attribute INIT_15 of inst : label is "899BBDDFEFE43FFFEBFCBFABF7FDFF6DFEDBDDFB5EED2A6FF5FAFD7E83DBC626";
    attribute INIT_16 of inst : label is "7BBF77BB4A9BFD6EBF5E76FD3A192064BC11C474A053442213A8A5A1C2380471";
    attribute INIT_17 of inst : label is "B7F7DFFFEDFEF77BBFD7E8382B8A645029A21509D452D0E11C02B88EBFE6DDDB";
    attribute INIT_18 of inst : label is "03D0F8BE0FC1C0F0F4F8FC7EF520152F88010E70D81C039FC46FBF7DEF4E38E3";
    attribute INIT_19 of inst : label is "7FFFF6FBD12CBEFE5FAAFB755DDDDFD1F378CEB2C9154578BB2D8C4DD9FCEE8F";
    attribute INIT_1A of inst : label is "6D777DBD7D87EF57EAF7FFDFF8E953D2FBFDACFF7D6FFEFBBF7B5BDFADFE8DF7";
    attribute INIT_1B of inst : label is "FBFD0A08FF3D8F3B24D9865E7F7FE9E28F4F40533BBDB6FCFB7FC8CDFD6FE0DF";
    attribute INIT_1C of inst : label is "BFFBBF8FF5F6FBD7BD1EF7BDEFCE7F739D87F8843F7DFFFDFC8FA57FB73A7F96";
    attribute INIT_1D of inst : label is "6FB2FBDEE1F877A6C9B7B2E19B97BE66E1D74F4FFA7A7E771CE3EE9D9D9CFDFD";
    attribute INIT_1E of inst : label is "7EF86233BFC7F3FFDE6E69931BC7D9C9AF5D78679F197F77BF3D243B7F34CEEF";
    attribute INIT_1F of inst : label is "4BDDDDDF9FABDE75AE5D737A7FEFDFCB74E5EF77EECFB5D5BBBD9DEDE1EFEEF8";
    attribute INIT_20 of inst : label is "FCFA4FD727DAA6587EBEA52C77D9EFEDF7D67CD5D7D44F77FFEA9D519C351E95";
    attribute INIT_21 of inst : label is "B8FD7F7DB66D3F277FDAFBFC7E077BFBDF5BE677CF6EF7DCFCB0EF866EF9FFB7";
    attribute INIT_22 of inst : label is "DFBF7EFDCFBF7EFDFB7FFEAFE844EEF7B9EF604FE6670F843BCFE447BF948B76";
    attribute INIT_23 of inst : label is "F7EFDFBF73EFDFBF7EFDFBF7EAEAA013F9FFFFF7F3FFF3FFFFEFEFEFEFE7F359";
    attribute INIT_24 of inst : label is "FEFEFEFE7FFE77EFDFBF7EE7DFBF7EFDFBD5D56FFFFFFF3FBFBFBFBF9FCEFDFB";
    attribute INIT_25 of inst : label is "F9ADFBF7EFC7F7F7F7F7F3FFF3BF7EFDFB9F7EFDFBF6AAABCFFFFFBFFFFFFCFE";
    attribute INIT_26 of inst : label is "CF9F575C7EFDF8FC6A7EFDFBF1F9FDF9FDF8FDF8EDDBB76EC7CF9F3E7CBABAF3";
    attribute INIT_27 of inst : label is "BF7FFF6FFB77EE44BDE03F7EFC7E353F7EFDF8FCFEFCFEFC7EFC76EDDBB1F3E7";
    attribute INIT_28 of inst : label is "E93589DF739DDDFE9E3BF8971DFFE6477F372AB3F7EFDADF7FF7DDEFDFBF7FEF";
    attribute INIT_29 of inst : label is "FEFF7ECF55DFB0434F9A73F79CBFFFDD7AA6FFEE7777FA7BFF9AC4F39DFFF5EF";
    attribute INIT_2A of inst : label is "BADFFD5FF33FFFEF3FFAFFFFFEEBFFDFDFBBEFEDDFFFF7FFD748FFFFE0697FF7";
    attribute INIT_2B of inst : label is "5BF8FFBF5FFBDFEBFFBDFEBAFEB9F7F5FE2FDA9FCFFBBF80662FB59FEF26FBC9";
    attribute INIT_2C of inst : label is "EFEF77FFEBEBEBE2DFDA6D9637EE1FC499307F9FC6FF7FAFFFFFFFFFFEE84DBE";
    attribute INIT_2D of inst : label is "FAB06A00FDCDFFFE9E1FFFECEFEF3FFFEBFF9FFFFF7DDC5BF8D3B873FF167FFD";
    attribute INIT_2E of inst : label is "3FFFF6DFDFB8B16EFEBFDE378F977B3ED6E7802BD305DF5FC7EF7E0AA9DFA7BC";
    attribute INIT_2F of inst : label is "DCBE57FBFA9B97CF7DEEEEF4925F7BEF5BB187BFB27E7CFFAEFBC810C5DE170F";
    attribute INIT_30 of inst : label is "FFFFB7F57D5F57D5F27BCEFBEB2FE13DDDBCFFFA3EF33D89BBF6CA7FFDFDFFBC";
    attribute INIT_31 of inst : label is "FFFAFE7BFFFFFF7FDFF7FFFAF4F1FF7FFFBBBF5E96FFFD7FFFFDFF37FFE07FFF";
    attribute INIT_32 of inst : label is "FFEF6EFFE7FFFBBBF9BFFF9F7FDD571DFFFFFFFFFBF1EFFFFF7F7FFF037FFE07";
    attribute INIT_33 of inst : label is "FFE7BFFBDFFEAABFEFFFFEFFFDDD8F7FFF57FFAAAFFBFFF5FFFD5578DFFFAFEF";
    attribute INIT_34 of inst : label is "FFABFEFF83FFD755EDFFFFFD6F21DFFFFFFFEAAB06FFFC1FFFF5DFF7FFFE7BBB";
    attribute INIT_35 of inst : label is "AAAFFFFFFF7FFFFFF7F7FFFFFFFEEEA5BFFFFFFFD774ADFFFFFD5540DFFFF9FF";
    attribute INIT_36 of inst : label is "FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA";
    attribute INIT_37 of inst : label is "B973FFFD7D70323FFD7BF59D4AC9C9AE7FF6BBE06BC9CAED6DD24B26783FFFFF";
    attribute INIT_38 of inst : label is "BADFACFDB6FF7DA2AEED6AFB5BBFAF6577E7BDBCBEB77BAD9BBFAEBEE84DF3FD";
    attribute INIT_39 of inst : label is "FF5D3FDAFFDC97DFB79C35FDEFD785DA5D7FEAF93F7FEFB6FD5D2CBAFFD7D7EE";
    attribute INIT_3A of inst : label is "3A2142814DB109D452D0E11EAEC05C29D29217DDF337CCDF33EDC274BDFCFF7B";
    attribute INIT_3B of inst : label is "9FFFBBDB69FF26A8F3FFF77D77FC6F7805EDFFB9FFCEE7FF0F4B9F9FFD6E8F20";
    attribute INIT_3C of inst : label is "0040CC80E048C982200F5F06FB7F30F2983E7CF9FBAEDFFF04BCDF79BAD1FF7E";
    attribute INIT_3D of inst : label is "0045100080002001404004040888004200000000007559001000000200011020";
    attribute INIT_3E of inst : label is "A0273807C8281E1100B0143FFFFFFDAD6BC5F40616B7577A0040400008000000";
    attribute INIT_3F of inst : label is "219FFEFEFFFEA19FFEFEFFFEBFCFFB7FF4728E01C8710E83024274000719507E";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "E837FBBF4A3A9428D7A74E6101999B9CD8CFB0410F2F0F7D46BE96EFDCEECBDA";
    attribute INIT_01 of inst : label is "F736EADD68F25AE6DC34F693DAC9B5CECE6CE557FE72AFFD3C9266EF7C4652FE";
    attribute INIT_02 of inst : label is "CBF3E5F9F2FDFEFDFBD4DB6DACDD493DEB335A4F3CE7C3B619A7192496DA66FD";
    attribute INIT_03 of inst : label is "F77F7BBDEB8636A699B9FC6F0D9AD28D9ACB71FDA9B2912E619AECE4FBDF97EF";
    attribute INIT_04 of inst : label is "C9ADAEE53BF9DF9AE734685E7FD9BD4571E71FF66B7F667B33FCC50DE6B3A277";
    attribute INIT_05 of inst : label is "D67BBA7DB9B7CFE90792D532BDDFAFE5BFEB12F5AAFBAEFAD7F7B7B7EF3F8FEA";
    attribute INIT_06 of inst : label is "F93D5899684A46A5A50FD6CB75FCF9E6EDF4081EFFF6CE4CE6EF656EE4980002";
    attribute INIT_07 of inst : label is "EF0D69558CF1AD2AB8EFA34ABBDBFDFDFF70F6A31B6F3F3F27DAB3279B5A3FC7";
    attribute INIT_08 of inst : label is "EE6FF0DA77AE7F1C3EB033235FDF697DF2E7F164F786B4AAFBAD4778D2ABA0E0";
    attribute INIT_09 of inst : label is "FFF7FC433FB6B8B17A1467D233FCD5AB19F7FFE873BFFCEDEDBDED62E7B387DA";
    attribute INIT_0A of inst : label is "F4FFFEE7CDBFE75DBFEA74DFF73FF777FEA7BA9FBB3FFFF7FFFF77F77FF777F7";
    attribute INIT_0B of inst : label is "FAE7E3D37FDCF9FFFD4EBEEF73EFFBDF4FB6F37FBFFFFEA7F4FFBEE7FDFFFEA7";
    attribute INIT_0C of inst : label is "FFBEFFFFFEFFEFBEFF9B53AFB3F73EFFFF53ABB3DCFBFEE9FD3FFFB9BFFDDF9F";
    attribute INIT_0D of inst : label is "FEFFFFFEFFEFFEFFFFFEDBFFFFFBFFFFFBFFFFFFFFFFFFFDB6FFEFBEFFFFFFFF";
    attribute INIT_0E of inst : label is "DF7DFFFF7DFFDFFDF7FBEFF7DF7DF7FFFFF7FFFFF7DFFDF7FF7FFFDDEFFEFBEF";
    attribute INIT_0F of inst : label is "EFBFFBEFBFFFEFFFFBFFFEFFFDFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFF6FB7";
    attribute INIT_10 of inst : label is "FCE3DFDFB2F9CE7FBE3FFD7FCA9D9EEB75F7BBED2ACFFFFFF7FFFDF7DFFDF7FF";
    attribute INIT_11 of inst : label is "F5A56F7ADEB593B5DCE8D9FB7304F01FC07E03F01FFC07E03BF01FEFE087BFB9";
    attribute INIT_12 of inst : label is "008FFFD59D7B6F1D4F3E91A257BFD36B6FAD65B3D9EEB77B2FF5C75FADF51DAE";
    attribute INIT_13 of inst : label is "5DFD6DDE436C7EEEDAFD3CADEBD6EBAFB8FBFC3EFA38CFBDFCF003CFBFF3F77E";
    attribute INIT_14 of inst : label is "FDEB26D6A967EA561825F7EB6EFDA9FA9F73B575F74034015E4DE20708421084";
    attribute INIT_15 of inst : label is "E34676B2DDEB64CDA754EBAD57358A3BA8737787BB55735DEEB77BBFAD4BB56D";
    attribute INIT_16 of inst : label is "6EF08ED55CD77BBDD6EAB2EF76C75EB7C37E1F7DCF9C7EFBF65F39CFF7C7DFAB";
    attribute INIT_17 of inst : label is "73B395DFDBBDDEEF77BBFB86FC3EFEE7CE3F7DFB2F9CE7FBE3EFD5AD3153BB0E";
    attribute INIT_18 of inst : label is "F03C0F83C0C23F0F0F0F878707E007F03FFB83FBFE23EFEFAD1DF3E6DA196596";
    attribute INIT_19 of inst : label is "EDB6D2326BD28A90E4EB4DF5BDDFF9AD0D4EFA873FC0180AF873775FF9AAF3F0";
    attribute INIT_1A of inst : label is "F4CD49B734B8ADBEEB186F5BEB3F187E1F0FCDD536DB416696F2CF528B2FBFA4";
    attribute INIT_1B of inst : label is "90FE07F074A1CA934F0930CEEE2E3F3EF1F9EFB6B6CE25959144FAAE44596AB4";
    attribute INIT_1C of inst : label is "2786B42C0607883882403DEB9C8AE09791B0D8E737216BE00060640968A0C594";
    attribute INIT_1D of inst : label is "48EC8FDAF4A50174496D53D55051954455305C5C12E2F6443FBFBAF5F2B398EA";
    attribute INIT_1E of inst : label is "49955591E0078602B5466946B21C09C952AACB5E52CF29AD6122644448C7A99F";
    attribute INIT_1F of inst : label is "5A54555E968B236B29EFB901DA95AF49AE8DBF24BBAF740427971CB9B1BFBB85";
    attribute INIT_20 of inst : label is "F1CAD6F8F4D762553E266B5CA4C7B7E136F9F3C5540B4D53FBFABFD49AAD7ABD";
    attribute INIT_21 of inst : label is "A6FCE7BF7B3978260087FF8D7D5E3976A0F20240C396E3CE2CCA4851017A0CFB";
    attribute INIT_22 of inst : label is "DFBF7EFDEFBF7EFDFA95150410636BDE759CFCBFA4A6A851E230A4B2242CCAD4";
    attribute INIT_23 of inst : label is "76EDDBB76BE7CF9F3E7CF9F155553993F9FBF7E7E3F7E3FFFFEFCFCFCFC7F35D";
    attribute INIT_24 of inst : label is "FEFEFEFE7FFF77EFDFBF7EF7DFBF7EFDFA8A2A0FFFFFFFBF3FBF3FBF1FAEDDBB";
    attribute INIT_25 of inst : label is "F1A9FFFFFFF7E7F7E7F7E3F7EBB76EDDBB5F3E7CF9F115404FFFFFBFFFFFFEFE";
    attribute INIT_26 of inst : label is "CF82A8A87EFDF8FE6B7EFDFBF5FDFDFDFDFCFFFEEDDFBF7EF7CFBF7EFD454413";
    attribute INIT_27 of inst : label is "B1A094CD28465FD97A663FFFFE7E353FFFFFFEFCFEFCFEFC7EFC76EFDBB1F3EF";
    attribute INIT_28 of inst : label is "DCFCD7AC88FDFF669DA33335D5AC8DF1E75541091B346D718545668D49DDEDBD";
    attribute INIT_29 of inst : label is "DE6F7FDE5FD8FB7C96E4EB1AC7BBE47C78F1D643F7FD9F67663E69C8F8D675C6";
    attribute INIT_2A of inst : label is "E91849BE6BB5D7CE69C6E6679B8C15151A9DBDBD8012401238BCECD8C893FBF6";
    attribute INIT_2B of inst : label is "5EFBBEF738A342898A34209F67D93EFCF93FFF1BE513372697E564F6ADFFAA7F";
    attribute INIT_2C of inst : label is "10E61FFFFFFFFFFF198C934964A2D5E7972FFBBDABDDEEF739FFFFFFEAABB3EE";
    attribute INIT_2D of inst : label is "FFFB7AD6FB4B70DEFDAD27B4B1D123DD8DA0909DFFFFFF63312EAB67667B6F1C";
    attribute INIT_2E of inst : label is "E592499A496285B5E274318C6A50C6A1B56C1B8813EDFF7B94F568A55CED260F";
    attribute INIT_2F of inst : label is "B589CD2A69B6B2F569A2597BE4CBFEAD332A57A627C9759464D6A74E34B552A9";
    attribute INIT_30 of inst : label is "FFFFC0A0A02A0A8287A5A90452179AFF136452F9A412E0A719FF996997956695";
    attribute INIT_31 of inst : label is "FF2FA99FFBFFFF7FDFFBFFFFF3FCCF7FFFFFF5F5FE7FFB87FDDFFFFBFFC07FFF";
    attribute INIT_32 of inst : label is "FFD5FA7FDFFFFB99FDBFFEFFFFFFEEFFFFF7FF7EFDFFE7FF80FFF77701BFFDFF";
    attribute INIT_33 of inst : label is "53E7BFF7FFFEBFFFE7FFB7FFFE1DDFBFFDAF7F9FEFFDFFEFFEFD56BF0FFF6BFF";
    attribute INIT_34 of inst : label is "C54A3FFEFFFFC57F7CFFF7FCB5796FFF3FFFEFFFFFFFFBFFEFF7EF7BFFD1FFFF";
    attribute INIT_35 of inst : label is "4150505FFBFFFF7EAF3BFFDFFDFFFFAA1FFEFFFDFFF754FFFFFC003FDFFF0FFF";
    attribute INIT_36 of inst : label is "F9F573FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEB741";
    attribute INIT_37 of inst : label is "D58B5FD395AB55B5FFADDB57BB1393316BFB4A334188CD7C92090A5651B778FB";
    attribute INIT_38 of inst : label is "D762B394DDF4375BB19B9B2CED6AB0DD8E5ED7D1C5CEE771B6C8B5C77BB7FB9F";
    attribute INIT_39 of inst : label is "5D632B1F7DBEBB6A9B5ABED6AD5B2EB0E79F4362E53E86EB15A6B1CF3E863ABB";
    attribute INIT_3A of inst : label is "C3FDF73E71FDFB2F9CE7FBE2B17BE03F3EFD5A88A1F287CA1FF395F7FFFAADF3";
    attribute INIT_3B of inst : label is "726B377FB3684706C6D64ED3BED7BEBB77FFFA9FAD5F2B5AEDAC1C5BFB8FB3FB";
    attribute INIT_3C of inst : label is "57AF559DF75F55FDCF7A085784040640032800BD2A088EFC5997F56FE9F5BEF3";
    attribute INIT_3D of inst : label is "FEEFBAFF6F5BFBFFEBEFFD7FBDFBD5FDFFDF7DF7DD820FB9FFE7AFDEFDFBBFFB";
    attribute INIT_3E of inst : label is "FDECFDEF3EEFB3F777CF778E7739CC314CFC06F7EFCF5ABDEAEB9FFD7BD5BDBF";
    attribute INIT_3F of inst : label is "F55288CB59AB755288CB59AB629969A2991F83F07C1F83E0EEF79EEFECFB7EE7";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "0200440CA35882145213B1ED50CCCDBE7E67E75DC212B643509256F9B001AAFC";
    attribute INIT_01 of inst : label is "FAEA76CAF46F2E5D4FA8BFDEFC2E20B8E5430916F1848DEF32D47F009264C451";
    attribute INIT_02 of inst : label is "2513329B89444A0685CFE787C72FB5C2F16EBD70BE1030090E53ECB64EB6DD7F";
    attribute INIT_03 of inst : label is "44C03C10F437AF75DCA574162FDDE82BDDB0FAC1DBC8DC5FF5DD1B7CD9CCCA6E";
    attribute INIT_04 of inst : label is "2FDF66419BE1BEC1F7BB854E6581D8293376270C260D7F6BFE01214EC1BF7138";
    attribute INIT_05 of inst : label is "1068305610810C0303097AAA1513BBB2C294D7B802EB2F4D3B137B00783C0A80";
    attribute INIT_06 of inst : label is "CB340EF697D56B7DFD853241248E8F3E9F37CCA9352269FFFF760C66ED40A8AA";
    attribute INIT_07 of inst : label is "260630E24660C61C4D264187026DB048610C1A80C403E3E3F6C02EE3D6BFB656";
    attribute INIT_08 of inst : label is "6914884FA32B308A0442D9B6844C3644C2B30E87130318710CC6393061C4424A";
    attribute INIT_09 of inst : label is "79977205980554B8174BB30A01864B7780A28A824BFF7EFEA12E10755AD82B09";
    attribute INIT_0A of inst : label is "D4B79DB769FC9579F63F7EFE4F285D7599B72E5A265A2515D4BD458EEC77665D";
    attribute INIT_0B of inst : label is "73768FBFC7AD9FFE366CB59E9B2D27B66FEC9B5FA637D937C4B3DD37C5B3DDB7";
    attribute INIT_0C of inst : label is "96D965B65965B6D9640CDBA574CFBFCFEED2BFD2F6EB4BADF52CF77FBCEFCADA";
    attribute INIT_0D of inst : label is "596C96D96D96D964965925A6D965A6D965B2496596596DB4926DA69A6DB6DB6D";
    attribute INIT_0E of inst : label is "EF3EFB4FB4D75EF9C73F9EBBDFFDFBDD74DB0DB4DB6CB0FFDFF1C73F965A69A6";
    attribute INIT_0F of inst : label is "B6D86597DF7DD75D7DF7DD75D6CF7CF7CF7CB7CF7CF7CF65B6DB6DB6DB6FFE1F";
    attribute INIT_10 of inst : label is "51B674725A9B5888D20488168B9CCA2D34D9CB1FD99FC9B6DB2CB2FBEFBAEBA9";
    attribute INIT_11 of inst : label is "841EDB97F57D79C37656A25FF350AFCB7731F95DC4B3F0DB8CAFC59D9B0CD15A";
    attribute INIT_12 of inst : label is "2A8946104EC5B9A9C7A3DD52405347F815BF22994CA2D249A65E05CA4AB0CFE4";
    attribute INIT_13 of inst : label is "465004930133E20A65C4226468D26986C0A734696E318C5338DFFC2AD8D2ADAA";
    attribute INIT_14 of inst : label is "C2B1684763BC60B448C42980249930DA29B24D36D83CC415185342F91CA739CA";
    attribute INIT_15 of inst : label is "8DB33F9A49002F3FE9BE94FE6DCDED19953E99F29F8C024924D149B6C1E9C402";
    attribute INIT_16 of inst : label is "733E67E3009249044A603A7DBA05C7AE45D435D2DCB6D3AE4B536B111A40B520";
    attribute INIT_17 of inst : label is "09C9F1DBE9245A29169B6C0BC071456E5B69E325A9B5888D205C109AFDA999A7";
    attribute INIT_18 of inst : label is "CEA7ACEB7ABE28ACA9ACD6D51C7FEC656CCD796E1BE05B4D84CE912FE74E32EB";
    attribute INIT_19 of inst : label is "16C97FFE600CBDB556579F9FD99BD7C5C6FCE5BB8C844006F8FBE0469AFC60AA";
    attribute INIT_1A of inst : label is "6373D58CC580D31D3F8DA5A01823F4471AA1DEAFEF2ED0FBFB3A69BA29268C56";
    attribute INIT_1B of inst : label is "69464604733101DA3234FBBC772F2393911D50016963D488EAD5005B3F48204F";
    attribute INIT_1C of inst : label is "9AF17B8A0C47851071100C6318DFC23E01BC717977454988400008CA988A6502";
    attribute INIT_1D of inst : label is "2696713DDA5FB526909621FFFBB5ABBABF972724193934933CE3CF0A98999554";
    attribute INIT_1E of inst : label is "B66FA805DC0301C15A68AFC109A39280E1C73BA56DE1DD12304008BB36024EC4";
    attribute INIT_1F of inst : label is "9FBEAFA905D1E377EC5FF213536566832C6FECB3ECFEFAE89A5CB26CC3EF6C7F";
    attribute INIT_20 of inst : label is "04B4397F791FE40FD3D81C62DB3B4B0C5174FFE8E6100224DEC13FE50FD0B530";
    attribute INIT_21 of inst : label is "B2F42383894D422600C8C025C20D7AEB10D9A415DFA2974C291FA7FFE4A0489B";
    attribute INIT_22 of inst : label is "D7FB5EBD7EBFDAF5EB8553AD9CF494611A462106C149F7FC19EAC9019851086E";
    attribute INIT_23 of inst : label is "FFFFFFFFF7FFFFFFFFFFFFFFBFFD500FFBFFFFF7F7FFF7FFFFEFEFEFEFFFBFDF";
    attribute INIT_24 of inst : label is "FEFEFEFEFFFEF5EBFFAF57EF5EBFFAF5FEDE5F4FFFFFFFFFBFBFBFBFFFDFFFFF";
    attribute INIT_25 of inst : label is "DFEDFFFFFFFFF7F7F7F7F7FFFFAF57FD7AFD7ABFEBD47F447FFFFFBFFFFFFFFE";
    attribute INIT_26 of inst : label is "FFE9E085FFFFFFF7FB7FFFFFFFFDFDFDFDFDFFFFEBD7FF5EBF5EBFFAF5BFFBBF";
    attribute INIT_27 of inst : label is "4FBEAF6E9BC62E40A000FFBFFFFBFDBFFFFFFFFEFEFEFEFEFFFEFFFFFFFBFFFF";
    attribute INIT_28 of inst : label is "793188E7A180C3BF8861984519E789833C514820F0E1CE4F2990FFEEBFF122B6";
    attribute INIT_29 of inst : label is "464A2A715A0D92EB225929B198D80BC89160C306030EFE3DB398C471872B867B";
    attribute INIT_2A of inst : label is "9ADC4DD7A16793042CBB5555586EA622DFFE26B272596C091830666C61612DA3";
    attribute INIT_2B of inst : label is "9960D33295FF9F77FFEBF7306C5A74F0E620982D40D798808D2B975FD2925EA0";
    attribute INIT_2C of inst : label is "040122AAA802A8060CD9619417AC314C0C180780C74BE5D2CE883FF575F52DB4";
    attribute INIT_2D of inst : label is "98802001A293A56EC2061B19382847226EC92422790140419AC2901C99101680";
    attribute INIT_2E of inst : label is "9B4D905CB296ADEAEEBD49D65DF52DDAF2CB002BD100E16EC446900AA37AA318";
    attribute INIT_2F of inst : label is "5CBA53171A09955E9DEE8AD4525529D35BE147D8F1322EAF2EEB7FF7ED5BF7F6";
    attribute INIT_30 of inst : label is "FF8048B7D8235D8A312DAA197DDB1418ECB14EB33725AB4CACC1CACF989A31A8";
    attribute INIT_31 of inst : label is "9FD7D19FB3F7FDBFE03F00D55AFA03B6FFFFEFFB6966F2BEFFFBF0DF64807FFF";
    attribute INIT_32 of inst : label is "FBF6933691FFFF7E867A9A03FFE858EEFAE7FFDFA96E764B3FFFF555FFD65807";
    attribute INIT_33 of inst : label is "AF99C3E0FFFF554396BB9FFFD85B71F11CAFFFD7F00432C0FFFFE807B71C74FF";
    attribute INIT_34 of inst : label is "FABEE72E07FFEAAA1E5FDFFEB50FFCB73FFFFAAAFFEE43FFBF141FFF3887FFFD";
    attribute INIT_35 of inst : label is "BBBBBBBD87FF7FFFF83F259FFFFAFAE7686CFBFFDDDEA65FFFFC003F30923BDF";
    attribute INIT_36 of inst : label is "CEBB9C0008CC6B902055B112888EE47A277B1B68CCEE44A375B912AFE6D54A3B";
    attribute INIT_37 of inst : label is "ED666E997F605166CDF8B8B5D7A185ACCDD236C040211E58D7CB4081102BC716";
    attribute INIT_38 of inst : label is "FBD1EAFFE66EA9977A4D76AE4A9F6A6BD7D5AEBABCDA691609277CD3EC2D56CC";
    attribute INIT_39 of inst : label is "7AD8631BE99817D7778837EA5CF707495377ABFCBFFDD5328F76AAA6EF7797CC";
    attribute INIT_3A of inst : label is "052B6B72DAB725A9B5888D21506C41E39190155450A146850BA980B418018C66";
    attribute INIT_3B of inst : label is "1F95E39320BB5120E36FD529F1EC0C1004CD3F21FE96C3BD18AA0C8249A68146";
    attribute INIT_3C of inst : label is "7FFDF7F3FD7DE7E3551B6300F2404812242840A0878AD66306AA4ED49A83363A";
    attribute INIT_3D of inst : label is "697CF7ADD4F5353777DF9F95DB9D1F731B30C30C336827DEB2FA7F7757CF7BFD";
    attribute INIT_3E of inst : label is "AAB6B7992B79582BED0ABC1A52B5A6F7E867FDA94659FE65DFF5E6D3DD2D5355";
    attribute INIT_3F of inst : label is "A115EEEA5FDEA115EEEA5FDEB668E7915012F04E3781F29C976CD7D516159502";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "E54AEF8DF713FDBB2B47467F93BA22C1F513F3EF842ECF75CABFF345FBBE3248";
    attribute INIT_01 of inst : label is "F713AAF569E2D3C675F52AF8AABC85DEEE6F8898FFC449F8B57A225F4ED781FB";
    attribute INIT_02 of inst : label is "FEFCFF7C7FBFBEEFBAD35D6EAAF4C7BD6B93DBEF2CF7D1F61CE55B6DB79B427D";
    attribute INIT_03 of inst : label is "F77D58A5697A129CF20DF5AF3C8AD2BC8ACB13ECA912F1F6278AEDA2FEF3FDF1";
    attribute INIT_04 of inst : label is "D9ADBDDD0D01093463FE6C5723EDBF2539F7BDF0686B225913B163ACD0B0EBB1";
    attribute INIT_05 of inst : label is "BFEFF403B0FAFBFED356D4F7EB7BBB6D2D7B38A57FFFFF5EDABDA2D6E96944CE";
    attribute INIT_06 of inst : label is "1CBEDFFD686B733F35C177DDEEAFADBFA9BE8FEBB687F97F44C5522774A8C00E";
    attribute INIT_07 of inst : label is "756DEADF255DBD5BEA75FB56F7DBEFF65BFD996DC55B2B2B2EEAD113A94A6AED";
    attribute INIT_08 of inst : label is "EE6B72263ABAAF754BE5F36BD0E9640E992AFDC63AB6F56F8AB5E3AED5BEE5FD";
    attribute INIT_09 of inst : label is "F7FF7D2956AAAB5FAB3C2AF7DD7C9D3A29F57D6D757FF15DF24CF324A595925F";
    attribute INIT_0A of inst : label is "BEFFBFB76FFFB759559B77FDDDB40FF7BFE5075FAF7FAFF77F77F777FFF7FFF6";
    attribute INIT_0B of inst : label is "FBB7EFFFF7FEE929A3CBFF3FF2FF87FDEDE6DB4BAE11FBF7FEFFFFF7FFFFFFF7";
    attribute INIT_0C of inst : label is "EFFFFFFFFFFFFFFFFB34BB656FFBB7EFF7B26546A48FE1DDFBBFFFCFB5F6FDDB";
    attribute INIT_0D of inst : label is "BEFF6DBFFBFFBFFFFFBFFFFFFEFBFFFEFBFDB6FBEFBEFFFDB6FFEFBEFFFFFFFF";
    attribute INIT_0E of inst : label is "DFFDF7DFFDFFDFFFFFFBEFFFFF7DF7FFFDF7FFFDF7DFFFD7DF7FFFFDEFBEFBEF";
    attribute INIT_0F of inst : label is "FFBFFFEFFFFBFFFEFFFFBFFFEFF7DF7DF7DF7DF7DF7DF7DFFFFFFFFFFFFBEFBF";
    attribute INIT_10 of inst : label is "45612728C00B18F6C03A344466BFA3F1FAB71AE5AFDFEB7DF7DF7DF7DF7DF7DF";
    attribute INIT_11 of inst : label is "132CE339C6338ABDC5F9AF8917EC6F107443A20D088744DE1F5F1231BE824543";
    attribute INIT_12 of inst : label is "0702C8CD5453AA2A5E3D51F5F897B52EB1F5E8F47ABD1F8FD5B54682E2C554BF";
    attribute INIT_13 of inst : label is "0FAD4FE35DD6C38BAF8795B972E77FC5A8057041340100C2E47FFF8063213DE0";
    attribute INIT_14 of inst : label is "696FA2D6B8B0FACC60C1B9AA7F0D417417F99FFAB571F24D7C1A00FC1886210C";
    attribute INIT_15 of inst : label is "5BDF52FC7E3FA4C933506B55373043E22EE4BEBDA9776CFE3D1F8FD5B07D934D";
    attribute INIT_16 of inst : label is "97D7AA5DDB3F8F47E3F51F6B63C6990D848000C6132C51051801631ED806E09A";
    attribute INIT_17 of inst : label is "FCBC882B0FC7A3D1F8FD5A89080315099628868C00B18F6C0370CDE5086621DC";
    attribute INIT_18 of inst : label is "3C0305C030BC1503000580041DBFFDA0055DF20CD9C3706F6F54E9D20E3DFFFF";
    attribute INIT_19 of inst : label is "CD36DB21530CCE92C5FD49EAB33A71071B431ED5766AB2AAFE627396BAAAF280";
    attribute INIT_1A of inst : label is "56C74EDC3EABED7CD53A7FDEEA2DF65B8D0D87D532DA42549FD7D5D45FD5ABAD";
    attribute INIT_1B of inst : label is "CE6544A6FEEE77FCA9A4A2CBDDFD2D2B0169123EB4822FEB93447EAC64FE2CB4";
    attribute INIT_1C of inst : label is "F587A645B1B16CE6CF6BDAD252CE92A4967364610A0A9D66BFBD03AD4BE6DF0B";
    attribute INIT_1D of inst : label is "BD4ADD9FF6F5BA4F066DC1B6CD9AD77736FBBF9FEDFCE81EFBFEDFAE3F7BD8EA";
    attribute INIT_1E of inst : label is "EDAD96C6B2FB76AEB1F03534BE5D40865CB3D7171887ADEDE44943FDEB7B3DD6";
    attribute INIT_1F of inst : label is "B8DDCCCC0215AFC93D4908AEA7F2550788DEFBBE776A774AF1DBEE5E7D5B5FCD";
    attribute INIT_20 of inst : label is "7BCDD6D3FCBA782D9AE5EB5EBCFFD3593ED3ED8BEBED84DAF6FB7BEE06EDFD7D";
    attribute INIT_21 of inst : label is "F4F7BAFD551FF9DFFFE77F9E7DF22D16EFEF7821C55C337FF87B7DDB3736A21E";
    attribute INIT_22 of inst : label is "DBB76EDDCF9F3E7CFB2BBEBEFC237DEFE97AFED68281BDDBE23582DE62A850F7";
    attribute INIT_23 of inst : label is "76EDDBB76BE7CF9F3E7CF9F3AAAAD953F8FDFBF7F3FFF3FFFFCFEFE7E7E7F359";
    attribute INIT_24 of inst : label is "FEFEFEFE7FFE77EFDBBF7EC7DFBF3EFDF9F5D5CFFFFFFF3FBFBFBFBF9FAEDDBB";
    attribute INIT_25 of inst : label is "F9ADFFFFFFE7F7F7F7F7F3FFF3B76EDDBB9F3E7CF9F6EAAAAFDFBF3F7EFDF8FE";
    attribute INIT_26 of inst : label is "CF9F55757FFFFCFE6B7FFFFFF9FDFDFDFDFCFFFCEFDBB76EC7DF9F3E7CAAFEA3";
    attribute INIT_27 of inst : label is "B16994386C2FD7D3BF0ABFFFFE7E353FFFFFFCFEFEFEFEFE7EFD76EFDBB5F3EF";
    attribute INIT_28 of inst : label is "D7F36FFB6F72B9466EDEEABF57DB766EC6279223AE5EB8BAF3C144D8898F2FE5";
    attribute INIT_29 of inst : label is "1EFD801E67F34516D5B6D66F45DFE4B76E9FFDBDCAE51DCA44F9B7EF72944E94";
    attribute INIT_2A of inst : label is "EC717F030C09FFD7F3DF6EEFBED9CF25B20967E5AD369AB696DF7BB7B2DE10D8";
    attribute INIT_2B of inst : label is "F6F69A3DF2CA4B29ACB6BAD6B5EAAF6F759FAFABBFBDCBA56BF5FEEEADEDBA7B";
    attribute INIT_2C of inst : label is "4A9D5FFFFFFFFFFDF74FDFBFBC4BC8EABF7DFFFD2CBE5F2FD600000FFFFFFB6E";
    attribute INIT_2D of inst : label is "FFFAF95523137EBF3CA6331116B44BF9D8C422CBFFFFFFBEEBB52F46444D5653";
    attribute INIT_2E of inst : label is "659361F2694BDEB56336B5AD6F5AD635A6E2AB27496FFFD377BF6F55F3AD1BE0";
    attribute INIT_2F of inst : label is "B7C8E57AECF6FAAD6F3378BFEDEBD7AD8E1AF7E604ED75DEF394EB7CA6B77BBC";
    attribute INIT_30 of inst : label is "FFFFA0888A208A222FB5FDB6DB133B5B13619935EAC0F5A7CEBC9C13F6BDAED7";
    attribute INIT_31 of inst : label is "EFAFAFFDFFFFFE7FD87BFFFFF5F5873FFFFFF7FD9E7FFF8FFFF7FFF3FFE07FFF";
    attribute INIT_32 of inst : label is "FBF7EEFFFF7FFEEE7BDFFFE7FF9EA7DCFFFFFBEEF7FFF7FFC0FFFAAAFF3FFFFF";
    attribute INIT_33 of inst : label is "D6FF9FFFFFFEAFF0E7FFF7FFB687EF3FFFDBFABFEE3BFFFFFFDD52AF0FFFD7FF";
    attribute INIT_34 of inst : label is "FFFFFE7FFFFFD556FEFFFFFFBFFCCFFFFFFFFD55077FFFFFF757FDFBFFF8FFFF";
    attribute INIT_35 of inst : label is "4451111FFFFFFF7FFFFBFFFFFFFDD7021FFFFFFFEBB20DFFF556AABFEFFF8EFF";
    attribute INIT_36 of inst : label is "B7777FFFFFFFFFFFFFFFFFFFFFFFFFFDFFFBFFF7FF8FFF1FFE2FFC5558EBF944";
    attribute INIT_37 of inst : label is "97189EF51D2D7489EBAB57571A3317E313D6BA32F412DE7284A641E78A9F7FAA";
    attribute INIT_38 of inst : label is "5762B3183D871B5DB3FB9B1DFD4CF3DD9E5AD4C1C7ABD1FAF6CCB7E35A92003E";
    attribute INIT_39 of inst : label is "9B46917D6FDEBB4A9316ECD5EBDAEEBCED934D62C610E36B15B7F1DB269E38FD";
    attribute INIT_3A of inst : label is "42D7084CB1828C00B18F6C01410483ED175532E8BB02EC0BB1A1E4F218044468";
    attribute INIT_3B of inst : label is "F26B1F7EB668265C8CC44476AE97EE52E3FA7ABBAD5DAB5A77A9EE7F7FC5A376";
    attribute INIT_3C of inst : label is "9E7B7FF379516F40749A025F8AAC68CB347FAFF5BB79EDFED5D7B74FECFC3571";
    attribute INIT_3D of inst : label is "616485A454153515575F9F15531D8B4102A08208232A054E803A3C2747844B35";
    attribute INIT_3E of inst : label is "4270067D015CC3DA9E08A81AC2358C691897FB8C6DAEAB8BD474A2929C295351";
    attribute INIT_3F of inst : label is "73F2BDD4ABAF33F2BDD4ABAF2CCB4D76561682804411024095081532B0ECD146";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "5451854015E77F9F1404C2E96844476A02203D75C57F99297001D32DDE4A4500";
    attribute INIT_01 of inst : label is "0F4390D0EC3E75CE33BC619D84CFB4C30F8AB08A1559442E2497080668061820";
    attribute INIT_02 of inst : label is "0307018380C164C9333438C861C2BDCEF984A7739EE3C43FEC5C9000969A4802";
    attribute INIT_03 of inst : label is "19B47831E500C05557D704090E21CA0E21D285521D12153681E17488011C060E";
    attribute INIT_04 of inst : label is "AB995A024CB5ADC8CE2DC3AD2F61603AE944C21A2D4613B09D96394B0075173D";
    attribute INIT_05 of inst : label is "852281C53E22070A841C2BA2118500474AD7B7AC0C73C665F3536C05CC98B418";
    attribute INIT_06 of inst : label is "1A0C18A3D1C4442961345C80422022203204F18448EC815577550846A64303F3";
    attribute INIT_07 of inst : label is "E80569520E80AD2A40E8A14AA26D200B8403D4E34304D4D4E0020442882940C8";
    attribute INIT_08 of inst : label is "8175F865F46643880444B78365D0EA5D00F40283740694A90CAD7F4052A4A0AA";
    attribute INIT_09 of inst : label is "99999C0320807C3815D3E4083A1C4B6683FD55603C00050213272037AA32049A";
    attribute INIT_0A of inst : label is "15001089524409C2444895200440A40944885220428001911919191911999998";
    attribute INIT_0B of inst : label is "04C8204020112200099301624480108910C964824B0040895100548950001489";
    attribute INIT_0C of inst : label is "1000040041001001017A4D8079544A020264C010993014A2544015324A09C220";
    attribute INIT_0D of inst : label is "0000900100100100000124100000100000000004000000000000000000000000";
    attribute INIT_0E of inst : label is "00800000800800020020000820000800000820800820000C0080002000000000";
    attribute INIT_0F of inst : label is "0041001001000040001000040008208208208208208208001041041041000044";
    attribute INIT_10 of inst : label is "167C02022DACA3538DC996A9941301A4C22505E1962000800820020020800824";
    attribute INIT_11 of inst : label is "027E52B5A56B6244400E1AA4621B62EC03941D10E4183B01E100E60401780125";
    attribute INIT_12 of inst : label is "C07E0B681314B2C1041FA04C301418869482C2603008040601691E28B4CC1048";
    attribute INIT_13 of inst : label is "B087190280D251B1A6A30073460F0601239947A643CEF50C03100238A92D0019";
    attribute INIT_14 of inst : label is "8AD73094DA9A5B61871B2638C80C16606200E0C0244EA04D01ACFD07E358D6B5";
    attribute INIT_15 of inst : label is "8ACF4829101926D9236B1FE2EB752C091112EA7CA4104210180D060120ED8219";
    attribute INIT_16 of inst : label is "5D4FA9041084061349841B62619E26D2BF45F1012CCF8A8845B5946A71BC91D0";
    attribute INIT_17 of inst : label is "D47661104203118CD462123E53D4049667C52822DACA3538DE45686FE498B022";
    attribute INIT_18 of inst : label is "C3E8F53C4F03FEFCFAF578F9E140015FC5D80D80001E4C304313C78843734734";
    attribute INIT_19 of inst : label is "CD36D264457A95D46610887C7321B3154CFBF5B41BD542A32E7B720824CC8E2F";
    attribute INIT_1A of inst : label is "33E2F58EF4685FA5F884EC3A76CA099460F0298BE8F648C57B898CA326B16794";
    attribute INIT_1B of inst : label is "F3AED7F2478199228D5E1C794D0DCAE01E5624E49D18D351CEEFB220AB3598EE";
    attribute INIT_1C of inst : label is "3BBE6E8E3C348BD0BEC01431087745AAE58CF3BDF9E87A1C006D392FD02984E2";
    attribute INIT_1D of inst : label is "2E63EE20213A75A2F13E78A9BA758AEEA93573501BCAC797155DD43DEEAAFBF3";
    attribute INIT_1E of inst : label is "79B24598280C6780EC2F9C820296DE71123ADDCCBEB919BE518870FC78F58518";
    attribute INIT_1F of inst : label is "6FBAAAB5C46FC25CD775F7289C39A8E0BDE75EF7759FBDB6BB7EBBDCB2547DE2";
    attribute INIT_20 of inst : label is "9DD3C81D257BA79261AB673A47891C37E91FD6B7980B66CA0A98D519E13C70DC";
    attribute INIT_21 of inst : label is "5CD6F440E9E48658FF1EC0E20304F8BF3F4BA73CF5235D600E148FA2E9C20CB8";
    attribute INIT_22 of inst : label is "244881027060C10206C5514113DE855A4E34C8BA38F04EA4A2B238B22F365BAE";
    attribute INIT_23 of inst : label is "8812244884183060818306095515241C0204080C040004080030181010180CA6";
    attribute INIT_24 of inst : label is "01010100810289122048910830608183048A0A30000000C0C040C040E0112244";
    attribute INIT_25 of inst : label is "0652000000180808080804080C48910204E0C182040C5550302040C081020701";
    attribute INIT_26 of inst : label is "3068A80180000303958102040E0202020201020710244881182060C10245415C";
    attribute INIT_27 of inst : label is "7CA68C2A298B18B24040C0000180CA40810207030103010280008910244A0C10";
    attribute INIT_28 of inst : label is "21E36E49B95304C9300228B91049AB82C89268A92B54A4F2CE28EFAA7DDDB7B6";
    attribute INIT_29 of inst : label is "385D800130114137D43EC229508024B32707B4C54C13206BEFF1B73959CCECCE";
    attribute INIT_2A of inst : label is "F89445C39042743824BA1110486F3886576F33B3C08240001BE1A8B0A0FA14D9";
    attribute INIT_2B of inst : label is "0D02A2822B75ADD617C85F25591458988308304C631706901CE2C76CDED9E692";
    attribute INIT_2C of inst : label is "00F707E00000000C114DFB9F27206928CB9464474F43A1D08EFFFFFC0002BED3";
    attribute INIT_2D of inst : label is "C008141150E099B186286C0E0FB1883EAF09C6BBE000010229F4A163EF456A1E";
    attribute INIT_2E of inst : label is "E7B365561BD8BC39B6358D635FB6717CD54B0243092500954666F9AF5A888C98";
    attribute INIT_2F of inst : label is "FB9CC197783F713AF9661C5C6DC5A55F1298862A93EC09A768BD1A95FDFA964F";
    attribute INIT_30 of inst : label is "FFFFE2A2828202000DA9AB248FCD2AEB15D634D08DFCCA6239025884C4CB3789";
    attribute INIT_31 of inst : label is "FFD2D67FFC0EFB7ADFFFFFFFF5F5FFFFFFFFEAAA97FFFFFFFF555F3FFFE06AAF";
    attribute INIT_32 of inst : label is "FAAF6FFFFFFFEEEFF9FFFF9F5FDFD71FFFF9FFFFEFF1FFFFFFBBBEEE03FFFF9F";
    attribute INIT_33 of inst : label is "D6E7FFFFFFFEAAFC7FFFFBFBF5D78FFFFFAFBFAFAFFFFFFFFFFFFD78FFFFFFFF";
    attribute INIT_34 of inst : label is "FFAB1FFFFFFFD7D5EFFFFFDD7F70FFFFC1BFBFFB07FFFC1FFF55F03FFFFFFFFB";
    attribute INIT_35 of inst : label is "5540001FFDFFDB7FE7FFFFE02FEFFE99FFFF01FFDFFD5FFFFFFD5540FFFFFF57";
    attribute INIT_36 of inst : label is "000000000C0038007000F001E807D40DAA1B5532AA05540AA805500004444215";
    attribute INIT_37 of inst : label is "8D7C249B2F5054C2479CB24F06B2972FB49A56C85A4BA1257B591198800A0000";
    attribute INIT_38 of inst : label is "0F6D7F27CBD9F6FF7DB7B7A74FD53DBBEEB9CCCDCB598CD43F117B1312DEA566";
    attribute INIT_39 of inst : label is "A4DF43806DBA3E45F70A1D98103C0E6AE1E3207DC9FB3EDB6BC6BDC3C667D9DF";
    attribute INIT_3A of inst : label is "FD5C24B33E0422DACA3538DEAF899C0AC803115C50F143C507218668E0050E05";
    attribute INIT_3B of inst : label is "3B676FACFEE980A69DDCC42E5E8C9100410793C71CE3CE79347A31CB46316C49";
    attribute INIT_3C of inst : label is "FEFFFFFFFFFFFFFFFF7FDF4392018A16C508003EE78A9E87158B3ED2F86E8628";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFF5D7FFFFFFFDFFFFBFFF7F";
    attribute INIT_3E of inst : label is "084BC188E2412D22657620F308E6118463380061BB47C5E5BFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "D0D182A21B1510D182A21B1526682EB410657EFFF3F27D1F64B568478BA24419";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
