-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu3 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu3 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "773081B9CD5EC954DD8919C57D5F5755555551CAA55555743171209B9B6A2EEC";
    attribute INIT_01 of inst : label is "2FBCAF556EEC53B341BB042B424AC136EC10AF2A9059C552351CAA5D0671548D";
    attribute INIT_02 of inst : label is "5EDA9412B9C01DB80B219550FCAEE56596955148D276EC1C56666F9F8242C661";
    attribute INIT_03 of inst : label is "88888888AAAAAAA88A8AA988BFFFFFFFFFFFA92316C3A9481269C5B0EA51049A";
    attribute INIT_04 of inst : label is "E6A4095757BC7A6A4B78D8DCF87BC7AE92F0948D7F09CE27104A494142000821";
    attribute INIT_05 of inst : label is "9DEE6372353FFF89FFCB9DEE60B2C124205EFB51489FA77E6A55655F9DC95277";
    attribute INIT_06 of inst : label is "A45221A210521013A0A153A05241F2B2627119A664A5DA609350557F0535C9ED";
    attribute INIT_07 of inst : label is "222202556477577474AA88AAAEEDFC07118A2492246582082EA7A6A5A4A7A6A5";
    attribute INIT_08 of inst : label is "4899D5550FB847371427044415718F3FB5CDD4F8C05103333012313103333020";
    attribute INIT_09 of inst : label is "2DF00C600D35C54D142A080AC1180C154765476562566765543350247F54BB49";
    attribute INIT_0A of inst : label is "00C02210E93030DCCD20C3CE88040E1C1023A303CF32C8CF7C903C043FF130F0";
    attribute INIT_0B of inst : label is "9E70106794C2794909DF00034000D0002C000B0001400070000C0008F30C300C";
    attribute INIT_0C of inst : label is "D7539F79A524275D496DA677D1719E70102794CE694909D75C77FEDE69D7D172";
    attribute INIT_0D of inst : label is "39E6029E554E419E516DD729A7D1729E5F59B49379F699D49DCD9750C9674909";
    attribute INIT_0E of inst : label is "989D0EEB4DFF779935DF7FEDAA72759D24275C6DC709A7D0729E42DD719A7D17";
    attribute INIT_0F of inst : label is "9DF41C2E5D28666D42A62D42A677D249DF6B2779B4DFF769935DF7FEDEA5D43B";
    attribute INIT_10 of inst : label is "99F04A9FA590755472A49E7195E69E6907579A49E5026008975026524275D5A9";
    attribute INIT_11 of inst : label is "79825275B499D56DC739A7D0729E5D43650949D4D77FFFDD25937926D14649C8";
    attribute INIT_12 of inst : label is "966DC719A7D1709E42DC739A7D0729E6039A524275B599DC6549E79A41D5A592";
    attribute INIT_13 of inst : label is "D07392639652427535DFFB79A4D955D532454D949493909D7519A6135DFFFF74";
    attribute INIT_14 of inst : label is "615736FDA964950D39A59D09D751965135DFFB49A6DD739A7D1729E42DC719A7";
    attribute INIT_15 of inst : label is "D28E598A4989D02255C199D098679837FFFED282690E5989D49D4D9D9D9D9DE2";
    attribute INIT_16 of inst : label is "7423556DE5DA426427196965DE709D4088948D855CDBF6A5945190269077FFFD";
    attribute INIT_17 of inst : label is "9D89D82E6571492641BD64B37FFCA4B249764B07B919074936FD9E4B0EFE2676";
    attribute INIT_18 of inst : label is "9279B64B07B9349F6ED9E4BFE2615736FDA9649DF7BFFFEEEECD2A49DFFFFD98";
    attribute INIT_19 of inst : label is "0000000111111111000008674DEFFFFBBBB34B92B7FFFF262762760B9D5D524A";
    attribute INIT_1A of inst : label is "44474E004CFB813BA78884B98799BB099958A88BC19B819958A8BC48A13B878C";
    attribute INIT_1B of inst : label is "0B1B8B0BA1002980320BA10010B1B8B0C00444474CDDC4774477445544554447";
    attribute INIT_1C of inst : label is "883BAA0B880B883BAA38883A9938BB38BB3A99388838880C00CC03BBA8BA1001";
    attribute INIT_1D of inst : label is "FD5CC5CFC45CFD5CF6CCCC4CEEC4CF4CEC44CEC4CD02BBBB23BAA2A884388838";
    attribute INIT_1E of inst : label is "000884402E6CC4DD5FFB473CF3CF3DD4DDCD5ECCE6CD6DCD56DCE6CC6CCCC4DF";
    attribute INIT_1F of inst : label is "883C880088AA88BB99B80012301133010B88B003F45200123019B45133012300";
    attribute INIT_20 of inst : label is "8070034E7400E77AC9778605C4AA4220FFFF00300003A1B819B2B33A288B88BB";
    attribute INIT_21 of inst : label is "C87C44E280784704800406B6E536140A50E14E4B8D47FC2B3DC35A871410D007";
    attribute INIT_22 of inst : label is "6CC8A2D480F0C270B492E0364B8D06288E87C62F24C462819206644CC6822C8C";
    attribute INIT_23 of inst : label is "7F28C47826828C426C9762C884E84E34880384070800E648ECF6C65CE4E4BF96";
    attribute INIT_24 of inst : label is "700066C0602ED262C1E62D1246C9A280006D9648E188442D8391B4E0C0088848";
    attribute INIT_25 of inst : label is "662685D468E24E368E668E8A6E2688226725D22362EAD6E2A66880E4E040A4A8";
    attribute INIT_26 of inst : label is "CFEDCFDCEDC00AAA47AA8B669680E1648E64E468421468024E468E426CEB26CE";
    attribute INIT_27 of inst : label is "888DA488E6523C79EB9E5A743D1982D110DC232730BEDFF155542020112FDCCD";
    attribute INIT_28 of inst : label is "2103210C4AA4F55557FFFFFFFFFFF9390089E77200B6776D822AE721ECC67CA4";
    attribute INIT_29 of inst : label is "2566559952495955565490555555552415554905514000506547654765476547";
    attribute INIT_2A of inst : label is "53C05C1A40171AA00500000146AEAABA9351AAA654D66A6A5AA5351699566949";
    attribute INIT_2B of inst : label is "0000000000000001650666515D999457AA05000105999058000016666505C501";
    attribute INIT_2C of inst : label is "EA940F94E43E94000055AAFF0055AAFFFAA5500FFAA5500016BC16BFE943E940";
    attribute INIT_2D of inst : label is "E94E4E38D2793940056F1B1B1B1B16BFA94E4E4E4E4F9500056BC6C1AF056AFF";
    attribute INIT_2E of inst : label is "8D379E49393A9500062222222C623F2DB2F888888889E50016C6D872CB1B1AFF";
    attribute INIT_2F of inst : label is "5B777924D3924DFFE2C61B1860889E4015ABC6C71C72D8722234EBFC0019B777";
    attribute INIT_30 of inst : label is "9630A426DA30ABC5B27788379BDDDDD5943D9DA390AC6B25B853F4B09CBE8094";
    attribute INIT_31 of inst : label is "00000003FFFFFFFC6C6C6C6C6C6C6C6FFFFFFFFFFFFFFFFF9393939393939391";
    attribute INIT_32 of inst : label is "C6559D555567B974BFF08B55FFF8000393939393939393939393939393939390";
    attribute INIT_33 of inst : label is "6DD75B75C61DB75CC51E17AD50B50BAF524333AF2BBD8594BC80BAB61C511752";
    attribute INIT_34 of inst : label is "93CB3E6F3C2EB3AEEEFB7A02E9EBF71A71979861F6DC75B71C5F75A7D97D861F";
    attribute INIT_35 of inst : label is "D716185D49F5F50043FEAB65F3F282820EBF9AE083F00FC226262626262625FA";
    attribute INIT_36 of inst : label is "D6003E2B95C410000810030C20810410000000800800400C20400C2058617527";
    attribute INIT_37 of inst : label is "79749D4D2713611585C7122041204F2C411B4520515050F2A5079050F6D5581F";
    attribute INIT_38 of inst : label is "81CD9149CF838F50F65974BE57F37A8251D07415241C1C163EBBB9271449C590";
    attribute INIT_39 of inst : label is "A07E5643E4646E7642E6649D554DD4541D75466951496E914A958081CE94EC80";
    attribute INIT_3A of inst : label is "F61D0712410791B4520539393B0CEC3014C2B004C1B00E6680B91A01E6680391";
    attribute INIT_3B of inst : label is "90AD2B31304D6F834008B041A919C955C71220412134520408C81EEEE07BBB81";
    attribute INIT_3C of inst : label is "C4C135BC84C4C119090FB05850F2E22C8185058FE22C81E1909A999C9C4C1190";
    attribute INIT_3D of inst : label is "81C870BE20701A05FFFFFFF8C5FFFA93E25D145B93E66145E846527E6A464243";
    attribute INIT_3E of inst : label is "424B90E3D4C7BECDEEC79E0E7E2AD79E8E8D53119092EAE53E8D5311937BEEC4";
    attribute INIT_3F of inst : label is "FFE4930C30450B82B8D34767252110545EE64DE251CEE2417BB241DC10263D4C";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "0011978741CE4F2C744F4741E338DF8BEC0EC8033FBEFB0040E3317871CCB9B8";
    attribute INIT_01 of inst : label is "1C542501400C023308EE0046A208CC1198013A8CF0072ED16C8033CC61CBB45B";
    attribute INIT_02 of inst : label is "760C99B7D36DB052DE97EC6C19D138F7205E30C48121B80BCF0F2A3A84C67394";
    attribute INIT_03 of inst : label is "333333330000000000000100155555555555D345BF9EC9914F916FE5B26453E4";
    attribute INIT_04 of inst : label is "033E8E377443C433C43CB4BA61C43C44F130764B4407413CC801F4F0C0000400";
    attribute INIT_05 of inst : label is "F453F6EB6C91545FFFC4F4D3F8F1401630131F8084F0B2C033CE487E4BC1E92C";
    attribute INIT_06 of inst : label is "BC8F8C7E8FBE9FAE4C4D8C4E8D8E5C4E6F8F173C041D73E0ECE100C08B0044DD";
    attribute INIT_07 of inst : label is "32100333300130213322301321123208F0F21B413C1E41000FBEBFBCBDBDBEBF";
    attribute INIT_08 of inst : label is "84FCB8C78AA62AA9AD8FA2000DCA469AA82AA0EA601233012012312023131021";
    attribute INIT_09 of inst : label is "1C70817F0C33E00C20F6281DC14C0C24675756446456564644554748C01C4F90";
    attribute INIT_0A of inst : label is "000002043FD0000C2BD0C30C22C3080F0C2350030C34084C30C01C2017381AC2";
    attribute INIT_0B of inst : label is "73E9709CFEEBDF974CBE000B0002C000B8002F000BC002C000BC0021030C2004";
    attribute INIT_0C of inst : label is "B8B171C77E5D32E2C5C7BD2C75C273E9709CFEE7DF974CB8B05FFD79DF5C75C2";
    attribute INIT_0D of inst : label is "273F8BFFE9CDE3FFEDD75C177C75C173E5DF5DF5CF1CF4BC4B06F8B47F92D78C";
    attribute INIT_0E of inst : label is "F24B8FDDE7FF5C5F5C79FFD717C12E4B5E32EDD75C077C75C273F975C077C75C";
    attribute INIT_0F of inst : label is "4BDC705FE7301BD7E57E97657F2C79ACB1E632CFDE7FF5E5F5C79FFD757E2D36";
    attribute INIT_10 of inst : label is "F3E02C3EDFF5C792A1BD73D75E9EF5DF5C7A7BD73F8DD20FF8B437E5D32E2E07";
    attribute INIT_11 of inst : label is "CF65D32E1FF4B9D75C277C75C273E2D1BE974CBA75FBBBA71EFDF7FE77A2A3C7";
    attribute INIT_12 of inst : label is "7BD75C077C75C073F975C377C75C373F82FBE5D32E1FF4B5D7B7BD77D71E9EF5";
    attribute INIT_13 of inst : label is "75C07FF2FBE5D32E9D7FF9E7BE5F9E2F1FF7C6F973767CCB8B3FBE79D7EEEE9F";
    attribute INIT_14 of inst : label is "E79CDF27E7BD73830797CB4CB8B0FBE79D7FF9C7BD75C377C75C373F975C377C";
    attribute INIT_15 of inst : label is "7309EF43CF24BA33C72074B27E3CF69FBBBA730DEF03CF2CB24B974BCB4BCBDF";
    attribute INIT_16 of inst : label is "2E9EEDE7FE7FE3FC3B7DE7BF7BC0E2D0C7FEFB9E737C9F9EF871763CFE5FBBBA";
    attribute INIT_17 of inst : label is "4B64B41BC7E1DB17E344F87F3BB8787D0F5F87D36F1765DF5F07E007AD6DFD2F";
    attribute INIT_18 of inst : label is "F9DF5F87D36F9DF5F17E0076DFE79CDF27E7BECB9CAAAA88889B13C676666DFE";
    attribute INIT_19 of inst : label is "00000000000000000008E5B2F72AAAA22226C4F19D999BBFB2DB2D06F1F876C5";
    attribute INIT_1A of inst : label is "74444E000671054004030401141111610151001055112501510005400440140F";
    attribute INIT_1B of inst : label is "54501454444444447754444445450144F0347444700134457445744574457444";
    attribute INIT_1C of inst : label is "14520751075107520753145314501450145314531453144F0074474775444444";
    attribute INIT_1D of inst : label is "20602612174320632720024133170272324503170E0011227520743314531453";
    attribute INIT_1E of inst : label is "5450147031702402402446402402403420024100170372024500173271301702";
    attribute INIT_1F of inst : label is "333D747602313120201274676474744541122773D55454545561156565767647";
    attribute INIT_20 of inst : label is "04706301006013120023040041332013557D6544444604015017356070310001";
    attribute INIT_21 of inst : label is "3140D41203204730060063200900D3309014012200720083220C3208304C1232";
    attribute INIT_22 of inst : label is "0324422324822324822224C3080030331047374314D11224D710504D2310504D";
    attribute INIT_23 of inst : label is "73000D3334054D3520D3160D20120132124C0063106013101033043013348323";
    attribute INIT_24 of inst : label is "70620106031053310D2200D212050106122093300D330049130D201C02312104";
    attribute INIT_25 of inst : label is "71333492001101620121013113234D720114D3340504D1013234D01402232034";
    attribute INIT_26 of inst : label is "021031031022321247100430902309020120133034D200610171015200137101";
    attribute INIT_27 of inst : label is "000C8000C8003210414415555155551555114444450010040002544567413131";
    attribute INIT_28 of inst : label is "7657464D5555E000000000000000057100B609FE00488BEBFEFBBEFFBBBFEBE0";
    attribute INIT_29 of inst : label is "1000000001000000000040000000001000002420050401406745745575667664";
    attribute INIT_2A of inst : label is "0006000002810000A081A4280000000001000000034200000000100000000004";
    attribute INIT_2B of inst : label is "00000000000000000810000A080002820060001800000A055556810000A08018";
    attribute INIT_2C of inst : label is "FFFFFAAA55400000000000005555555555555550000000000001555555540000";
    attribute INIT_2D of inst : label is "FFFAA540FE954000000055AAFF00555555500FFAA55000000000156AAAFFFFFF";
    attribute INIT_2E of inst : label is "FA940FFA95400000005AF05AFC03EAFC05550FA50FA5000000156BF015AAFFFF";
    attribute INIT_2F of inst : label is "005AF1AC1AC5BC0003A4394F94FA50000000156AFC056BF05AF16FFC0390E943";
    attribute INIT_30 of inst : label is "1DF0E2404DF0E19005AF1694000FA5001B06A505B0E539400776215A50888900";
    attribute INIT_31 of inst : label is "FFFFFFFFFFFFFFFC0156ABFC0156ABFFFFFFFFFFFFFFFFFFFEA95403FEA95400";
    attribute INIT_32 of inst : label is "C2EA6AE009B24E807FC0C755555C0003FEA95403FEA95403FEA95403FEA95403";
    attribute INIT_33 of inst : label is "27F309FCF38A9FC2E10A4B4FB4BD2F68E19180768EF4AE907F52F69E4F233301";
    attribute INIT_34 of inst : label is "C80CB4378131889393D3B4CBDAD3AF4AF09F49E4C27E309F8F2AF8AF09F89E4C";
    attribute INIT_35 of inst : label is "AECA792D04ABB000A29787A7E2912163A7B46FD082F00EC2A2A2A2A2A2A2A2D0";
    attribute INIT_36 of inst : label is "023A013855C01002041040000000000000002041000082041041000029E4B412";
    attribute INIT_37 of inst : label is "F0333F0CCF8323DDF00E21100038281010330050332008013593C02C15E024C0";
    attribute INIT_38 of inst : label is "5441BB464E2A63D8800EF07D578BF12580A023351B73733A00C44EFF423FD08C";
    attribute INIT_39 of inst : label is "05402050020540105001054010500105000054001F9104447D34755440994475";
    attribute INIT_3A of inst : label is "580A22315803C330050295402F90BE4511000501080520101440405100014400";
    attribute INIT_3B of inst : label is "702B9EE0A0171B4A87347000478787330E211000333001028F140DDDD0377740";
    attribute INIT_3C of inst : label is "82805C7F76828057978F6C70F803D13840C74F81D13840F57574787878280579";
    attribute INIT_3D of inst : label is "C0E2605F500801C35555555E8C0003600D744003600DD4003CD5F5D1F1E1F1C0";
    attribute INIT_3E of inst : label is "C1D7781BF6DF460761F37D8DD215D37D856FDB30707111DD066FDB3071C861F0";
    attribute INIT_3F of inst : label is "5555030C30A80E43A4B2293D3F94A6E2AFD3C7D3C78FD3C7BF53C7C00C39BF6D";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "19A8CD0D23448D30D84D4D63549F260C70E7062335C71C18021830D0D34CA032";
    attribute INIT_01 of inst : label is "14813408955A8AE86604880C592BA1992220218CD48017080462334ED005C201";
    attribute INIT_02 of inst : label is "84121658555255952159518DBAC992545824920E23983227267E79F9E3E3FB42";
    attribute INIT_03 of inst : label is "0000000000000000000000008000000000001515552521629556554A4858A555";
    attribute INIT_04 of inst : label is "433CDF9890410433CEC0101603C41048F380D641840D2234E403E262D0EE4100";
    attribute INIT_05 of inst : label is "DC23704B0570008D4038DC235AC002133CAB8C458891304433EE04B2C1234B04";
    attribute INIT_06 of inst : label is "092B3B39382B0A0929282B2A29283B2A1904033C803CF3C9F25062449506D028";
    attribute INIT_07 of inst : label is "3012330120123120131310203210330040E336211434F80F37090B0A080A080A";
    attribute INIT_08 of inst : label is "889812DBB4C2F4C35CCA6F042EF5F824CDDA93C2B09333000111122333001223";
    attribute INIT_09 of inst : label is "F0421015C00200010600001F0009B00103322111310201102023300395642045";
    attribute INIT_0A of inst : label is "00000005014C00011D4C00000000000C0043004C308008B00002000200307100";
    attribute INIT_0B of inst : label is "5344D704D2334D0C28130000C00030000800010000C00030000C00000C204000";
    attribute INIT_0C of inst : label is "108093413430A042034D3704D34C5344D704D2334D0C2810823554D14D34D34C";
    attribute INIT_0D of inst : label is "C535ACD3434348D3434D34D534D34D53435D35D35D35D8168128D0828D204C28";
    attribute INIT_0E of inst : label is "DD81E3234D55741D75D3555D077A048130A0434D34D134D34C1354D34D534D34";
    attribute INIT_0F of inst : label is "C135D3034D33034DB1344D303504D5141350904D34D55745D75D3555D1742088";
    attribute INIT_10 of inst : label is "56A04F6A14534D02C004924D3514524934D4514926434C8CD08233430A04200D";
    attribute INIT_11 of inst : label is "49930A0434DC134D34C134D34C13420A364C2810D373330D54D34534D2C72684";
    attribute INIT_12 of inst : label is "534D34D134D34D5354D34C134D34C135ACD3430A0434DC134D4514924D351452";
    attribute INIT_13 of inst : label is "D34C135CD3430A0434D55345348D3422A34D28D0C0D0D281080D34D34DCCCC34";
    attribute INIT_14 of inst : label is "4D36378DC924C9D90D4981281081D34D34D5535534D34C534D34C5354D34C134";
    attribute INIT_15 of inst : label is "D3355DB75DA41E375D11D810D375D5373331D3355DF75DA012811D8141410123";
    attribute INIT_16 of inst : label is "04B0434D34D34334B0D34924D359C20BF8DEC134D8DE372491D0D375D1373331";
    attribute INIT_17 of inst : label is "411412235DC748155D274001B333B0088D7700188D0D135D378DC0806E8E3605";
    attribute INIT_18 of inst : label is "54517700188D35D378DC0808E34D36378DC9244174F3332222000449D88888D9";
    attribute INIT_19 of inst : label is "048C048C048C048C08E500105D3CCCC8888001127622223640440488D771D205";
    attribute INIT_1A of inst : label is "12221C201202122212211222121221222121111211212221211121121222121C";
    attribute INIT_1B of inst : label is "12221212121212120112121221222121C2121222122212221222122212221222";
    attribute INIT_1C of inst : label is "12111111111111111111121112121212121112111211121C2111202011212122";
    attribute INIT_1D of inst : label is "10100101010110110102002011010010102021011C2111101111111112111211";
    attribute INIT_1E of inst : label is "1111110210120220220200200200220202002022010010202022011010100101";
    attribute INIT_1F of inst : label is "103C101020101010101010010202021212120103D11111111111111111111121";
    attribute INIT_20 of inst : label is "50406106406067A400B5000000444744003D2121212112212211011111112121";
    attribute INIT_21 of inst : label is "76E000094B6504140690635810610351006C06BA00EA6007E900F700F00009B6";
    attribute INIT_22 of inst : label is "A94003614003614003614003004094B658047EE5D00BED910E6ED8007E6ED500";
    attribute INIT_23 of inst : label is "47E600F7EE6D00FED10BED005065067254005061406065006B9800B7A9800B7A";
    attribute INIT_24 of inst : label is "4061180631810B1110B111033910540675810759107668107510506009B765C0";
    attribute INIT_25 of inst : label is "F21C8100C06006C00690067BE5DC00EEE9D10FEEED910F7E5DC00064094B6640";
    attribute INIT_26 of inst : label is "544477766659B764047604E10FA810D006006BAA810D906006D006D00069C006";
    attribute INIT_27 of inst : label is "5550055500154000000000000000000000000000000000000000647654476655";
    attribute INIT_28 of inst : label is "7657766155550000015555555555554200000130000013000000000000000005";
    attribute INIT_29 of inst : label is "2005AA50058401555401600000000058C000042001C800625447665477654765";
    attribute INIT_2A of inst : label is "23C185A5A440A9AD18D55544206DBE7905039394006106FF0E4058006BFE9016";
    attribute INIT_2B of inst : label is "0000000000000000042E94018BA50042001C80062016B104000063E94010AF87";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "5555555500000000000000000055555555555000000000000000000000000000";
    attribute INIT_2E of inst : label is "55555000000000000000055556A95556AAAAA555500000000000000555555555";
    attribute INIT_2F of inst : label is "00000556AABFFC0003FFEAA555000000000000000155555AAAAFFFFC03FFAAA9";
    attribute INIT_30 of inst : label is "015A540016AFA9000000555555500000005555555A554000005AF00000FA5000";
    attribute INIT_31 of inst : label is "FFFFFFFD55555554000000015555555555555555555555555555555400000000";
    attribute INIT_32 of inst : label is "891951CC69666578501DF8930002AAA95555555400000003FFFFFFFEAAAAAAAB";
    attribute INIT_33 of inst : label is "9C9667258A807261988192394E60BE350332C8B08EE2514853AFE371988E3213";
    attribute INIT_34 of inst : label is "E62EE33268BA63D9998E23CF8C8E42672262651999C966725884267226265199";
    attribute INIT_35 of inst : label is "61D146498218440036784214E670193B387C0764C17405D1999999999999988C";
    attribute INIT_36 of inst : label is "58C764B424001040000004004008300108081041041000000000000005192E08";
    attribute INIT_37 of inst : label is "26658899622678521EE3538C890EF23012E311B4A8022D937802548DB0818905";
    attribute INIT_38 of inst : label is "691D15185C201A881D6D48529F1AA010348225044105050365E26462E7589994";
    attribute INIT_39 of inst : label is "1101C190141101C190141101C190141101C190504550754191519A691E16519A";
    attribute INIT_3A of inst : label is "034812E000466E311B4800001145451100701900501101C0640501101C064050";
    attribute INIT_3B of inst : label is "D031CF7BC00D0F5BDBA120424D4D4D69E3538C890E31134BEFAD2F7F70BDFDF2";
    attribute INIT_3C of inst : label is "EF003400B5EF004D4D347A7E3DAB844D62A7E3DB844D62D8D8D4D0D4DEF004D4";
    attribute INIT_3D of inst : label is "32927637008721890000000DA056A4F5931465A4F65344523623435353535340";
    attribute INIT_3E of inst : label is "336D0975C250DD4DD0650FD435F0750F9BD40980D0DFB0425DD40980D355D064";
    attribute INIT_3F of inst : label is "002AA91ED1078FE3D0134737347915444FE34D134D23234D0CB34D40203F5C25";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "5024030300D3874C70C70300C7F1FFD30D80D8031C30C35174CB003031C01EED";
    attribute INIT_01 of inst : label is "04C20C0FC009042410BB417704109042ED05DC0C781700C13D8031D485C0304F";
    attribute INIT_02 of inst : label is "003C0000000003400000033C1C111FCBF03FF4C10073FD01FD81850510104D04";
    attribute INIT_03 of inst : label is "4444444444444444444444447FFFFFFFFFFF003C00000000000C000000000003";
    attribute INIT_04 of inst : label is "331C0DFFFD36D331E07CF8F070D36D387030304FD303031D0000D0D0D4500000";
    attribute INIT_05 of inst : label is "7631E3C13C1800C7403C7631C3DBB0707831171C0074D3D331FFD8FF8F00C13D";
    attribute INIT_06 of inst : label is "5477675777464646464675457565445474DBCB1D300C71C0D0C03FD383034E30";
    attribute INIT_07 of inst : label is "2333330001111223330012233012230DBCD001001C0FC3C20857565656555554";
    attribute INIT_08 of inst : label is "007CFFFFC33093330C1E09000FF0C3E337CCC030903000111111111111222222";
    attribute INIT_09 of inst : label is "C0411010C00202200000104F002D700776666665475464445477577EC0FC0718";
    attribute INIT_0A of inst : label is "03000001000C0001080C00202200004C0003040C008008700002000200305008";
    attribute INIT_0B of inst : label is "B1C0302C7002C7D704F70001800050001800040001800050001C00000C104030";
    attribute INIT_0C of inst : label is "FDBCB1CB1F5C13F6F0C71F3C70C0B1C0302C7002C7D704FDB01C0072C70C70C0";
    attribute INIT_0D of inst : label is "0B1C00B1F0C0C0B1F0C70C0B1C70C0B1F1C71C71C71C7CF04F487DB087E3D704";
    attribute INIT_0E of inst : label is "70CF0331C7001CC71C71C00731C13F8F5C13F0C70C0B1C70C0B1C070C0B1C70C";
    attribute INIT_0F of inst : label is "CF1C3031C70031C7C31C07031E3C730CF1CC13C71C7001CC71C71C00731F6C0C";
    attribute INIT_10 of inst : label is "77B0177B1C71C700701C71C71C1C71C71C7071C71D00C00C7DB031F5C13F6F03";
    attribute INIT_11 of inst : label is "C705C13F1C7CF0C70C0B1C70C0B1F6C21C1704FC71CCCCC72C71CB1C775B0780";
    attribute INIT_12 of inst : label is "B1C70C0B1C70C0B1C070C0B1C70C0B1C00B1F5C13F1C7CF1C7071C71C71C1C71";
    attribute INIT_13 of inst : label is "70C0B1C0B1F5C13F1C7001CB1F870F6F21C3087D7030304FDBCB1C31C733331C";
    attribute INIT_14 of inst : label is "C71C1D07471D7FC3030FCF44FDBCB1C31C7001CB1C70C0B1C70C0B1C070C0B1C";
    attribute INIT_15 of inst : label is "7002C702C704F031C30038F0302C701CCCCC7002C702C704F44FC78F8F8F8F31";
    attribute INIT_16 of inst : label is "3C13F0C71C71F31FBC71C71C71C2F6C3FC704F1C70741D1C7C30302C701CCCCC";
    attribute INIT_17 of inst : label is "8F0CF071C731D301C741D0170CCFD014071D0170C70301C71D0747010F331F3F";
    attribute INIT_18 of inst : label is "71C71D0170C71C71D074701331C71C1D07471F4F1E4CCCCCCCD701C073333470";
    attribute INIT_19 of inst : label is "0888CCCC00004444A50000E3C79333333335C0701CCCCD1C23C33C1C71CC74C0";
    attribute INIT_1A of inst : label is "01012E200101010001000100010100100010000010101000100001010100012E";
    attribute INIT_1B of inst : label is "01000101010101010101010100100012E2010101010101010101010101010101";
    attribute INIT_1C of inst : label is "01000100010001000100010001000100010001000100012E2010101010101010";
    attribute INIT_1D of inst : label is "00100101010100100101001010010010101010012E2010101000101001000100";
    attribute INIT_1E of inst : label is "0101012200100100100100100100100101001010010010101010010010100101";
    attribute INIT_1F of inst : label is "123C100010101010101010010101010101010123C10101010101010101010101";
    attribute INIT_20 of inst : label is "00002402402020000000000000645765FFFC1010101001001001010010101010";
    attribute INIT_21 of inst : label is "0040000514000044020024400240244020200200000000000000000000000540";
    attribute INIT_22 of inst : label is "0000040400040400040400040000514000000440400044002444400004044000";
    attribute INIT_23 of inst : label is "0040000044040004402044004024024440004024402024402000000000000000";
    attribute INIT_24 of inst : label is "0024400244002044020440244002440244002440024440024402402005400000";
    attribute INIT_25 of inst : label is "0440002400240204020402004040004040402040440020040400002005140000";
    attribute INIT_26 of inst : label is "7777666666654000000000002000020402402000002000240204020440200402";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000554444477777";
    attribute INIT_28 of inst : label is "7776666000000000000000000000000000000030000003000000000000000000";
    attribute INIT_29 of inst : label is "30000000018C000000005300000000108000042001C800727776666655555444";
    attribute INIT_2A of inst : label is "2411480000520000104505041001554001C55400005000005000100000000007";
    attribute INIT_2B of inst : label is "0000000000000003C52AAAA109555442001C0007200001CC0000620000188005";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000155540000000000000000000000000000000000000154000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000055555000000";
    attribute INIT_31 of inst : label is "FFFFFFFC00000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "415DD97FFF5344501001FDFFFFF1555555555555555555540000000000000003";
    attribute INIT_33 of inst : label is "1B5106D4401F6D40501DCD097C6C0D06F0CE40D40C505C6013C0D06DC43B1100";
    attribute INIT_34 of inst : label is "3008500700220E51D142D03343426D47D07D47DC41B5106D4436D47D07D47DC4";
    attribute INIT_35 of inst : label is "5D0DF70400D74000F01202DF3017070702003338001800619999999999999B40";
    attribute INIT_36 of inst : label is "3C0300203F000000000004004004000100000000000000000000000037DC1003";
    attribute INIT_37 of inst : label is "D0C1343C4D0E304C14C30004004C900038B3380E30C03C001F014C3C10BFFC30";
    attribute INIT_38 of inst : label is "0038003BCF0701C1CCF45013FFC1E000F3C03D7F0D71717F0044474D0D134345";
    attribute INIT_39 of inst : label is "380343403434030300303003C3C03C3C038380E0E000D003400300003C0003C0";
    attribute INIT_3A of inst : label is "FF3C03B0C0C14B3380E00000000D003400C03000C03003C0F00F03C0380E00E0";
    attribute INIT_3B of inst : label is "30DF0D3240073702C3082000030303F3C30004004B1300C33D038CC88C332220";
    attribute INIT_3C of inst : label is "C9001CC0D0C9000303C4DC0C0C02300410C0C0C1300410C0303030303C900030";
    attribute INIT_3D of inst : label is "20C030D80C020043FFFFFFFCC300013004C0E38130040E3807C0C0C0C0C0C0C3";
    attribute INIT_3E of inst : label is "F0F1FC31B06C04074071FCC7D0C071FCCCC7C1B03C3CC07F04C7C1B031C04070";
    attribute INIT_3F of inst : label is "FFFFFFFAAACF0DC344F10D1D1C103020F331C731C30331C3CCD1C34F03371B06";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
