-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FE7FCF84164E499F999D1A4BE59C93909F8BE8FE07F3BEBC9F958FE737CB6765";
    attribute INIT_01 of inst : label is "8F30549FFAF3BA6430975FFDF364F322FECEDF25737F2762FFB39C9D8FB9CC39";
    attribute INIT_02 of inst : label is "00D588187F6140AF84123F51A523FD3B44A32324967FB49970FBEC80A0D33B00";
    attribute INIT_03 of inst : label is "B8712C13DF73F4FBF3E3F2B92F9F9CCECDD64DA739FA99FF5CA8BF57D5F42088";
    attribute INIT_04 of inst : label is "7FD7E59EED5AE2D4B797AAABFFFBFC100904027F19375939279EBEBFB9CB5879";
    attribute INIT_05 of inst : label is "DF43EFEF777AC077189E7FF3F67FD977EE3FBFCFBA6FD07F1BE43F0DFF9DDABD";
    attribute INIT_06 of inst : label is "17FE4119C3021900964DC8232823249A37239044C9B552120BA7FFFB53FE588F";
    attribute INIT_07 of inst : label is "0C51624FA03E124924924924524FA003081187FCDB7F9E30C9F1FD6494B23FAC";
    attribute INIT_08 of inst : label is "FA80AA8D400051ABAFF451080D222828BE8A51408111DDFF6CB3CFFEAE3E7499";
    attribute INIT_09 of inst : label is "D9667E2BFFEF7293FFD20C0DCD3C5FFE09FED98D22DA5E3DA5E20D2452D22DAF";
    attribute INIT_0A of inst : label is "42B7C0822010A75555C8848A867D02A58EAEBF9FF9F7FB3FB33313F1BE02D37C";
    attribute INIT_0B of inst : label is "965F70FFFB2CFEBE7FE23E2C8896254D5F3FDC2F1CF88E7AC2B85FA100423ADC";
    attribute INIT_0C of inst : label is "DE6DF7EBB3C537DDF5CBBA6F8EA2F9A8A89DC6E935337DB8BFFFE09A90FFCF39";
    attribute INIT_0D of inst : label is "23C1A6F9B2934544EE3749AE6BEEC5FFFE3BC2C91A0D31623CC2CE907989E399";
    attribute INIT_0E of inst : label is "8B8B89FEA166359A79A3FA49A1FBC66D6687C78133270C626031D23196460FC1";
    attribute INIT_0F of inst : label is "00000247F2000000AEEDE016AA60880A0000016AA8F66667E758EAAEF759FFF6";
    attribute INIT_10 of inst : label is "BF3566D2B8FC000000000000000731200000026CA042FC436484C6C90E1CC480";
    attribute INIT_11 of inst : label is "1B91AFE3215FFDF13F8E0053937EB3EB3C9733C01FDCCE1BF2499B930E39717C";
    attribute INIT_12 of inst : label is "AAA80554000C03DF09E53815C29C72BC9FD64D53AF57B1C10B0000057A9C10B3";
    attribute INIT_13 of inst : label is "D3B4ED3B4ED3B4ED3B4ED3C02843FFFFEFAABFFFFFFFEAAAAAFFE6AAABFFEAAA";
    attribute INIT_14 of inst : label is "219861FB002440B002C00B4ED3B4ED3B4ED3B4ED3B4ED3B4ED3B4ED3B4ED3B4E";
    attribute INIT_15 of inst : label is "FFBFFC77DC4183FC4183FC10180FFC10180FF9DD18F87F2187F1060FF08181FF";
    attribute INIT_16 of inst : label is "CC27FFF0C5FFF799EFC87984DF6EBAD9B7E78DD2E0FD5949F3F011AAFE96EB7C";
    attribute INIT_17 of inst : label is "4B335AD430E60E41A40F0800C00E41A50060006FDAE8F913E11A5F800000800F";
    attribute INIT_18 of inst : label is "3F3D8BBFFB999FF8E471FFBCFC18A338D7FCC38DFFFD2C973CDFCDFA542FECEB";
    attribute INIT_19 of inst : label is "81AEB556001733202EE3929285DC9FA4FACBBCFFFB21196785C5FB27F87F63E5";
    attribute INIT_1A of inst : label is "DB94FBD6DDDDDCDC5DC6A6CCDE532AAAAAA3AFFBAF91E78099C4FEFBFE878E53";
    attribute INIT_1B of inst : label is "55C2B33B7266DF2D6657A44FF3EFB719661EAB7A6FAAAAAABA80F7CDF5CFADCE";
    attribute INIT_1C of inst : label is "E3DC7CF8F71F8AF57B87DEAF71FBD5EE1F7ABDC7EFCF71F3FEEAFEAAC9BBEEEC";
    attribute INIT_1D of inst : label is "FFD7972FBC03060DEE5E1FAAFB979F55EE5F78F73FBCA7B979EABDCFCF57B97D";
    attribute INIT_1E of inst : label is "DFFBBE9FEDDF7FEBCB8FDEFFDDF4FF6EFBFF5EDC3EFDF4FF6EFBFF5E5C3EFBBE";
    attribute INIT_1F of inst : label is "DF7FEBCB9FDFFFDDF7FEEFA7FB77DFFAF2E7F7F77DFFBBE9FEDDF7FEBCB9FDF7";
    attribute INIT_20 of inst : label is "F4FF6EFBFF5E5C3EFBFFFFFDDF7FEEFA7FB77DFFAF2E3F7FFFFF77DFFBBE9FED";
    attribute INIT_21 of inst : label is "5FDF1515FFACB24B368001F83F00014003F00107C18F73F8AFF7FFFFFBBEFFDD";
    attribute INIT_22 of inst : label is "69C45F20F136E269DC05B4FBA99BF9B267F20E044CA77C7FEC448BEBFE722CF8";
    attribute INIT_23 of inst : label is "96665570000019C447DC2B3FC64C415114326D3FF50DFFC474EBF47F2283E42D";
    attribute INIT_24 of inst : label is "C4BF5A28AFA625FAD3457D312FD68A2BE9897EB4D15F6E258962589625896258";
    attribute INIT_25 of inst : label is "12C760080FB8567E8C988C9FC7479FE4759D55C00FEF4554BA977897EB5D15F4";
    attribute INIT_26 of inst : label is "5FF0D02D2BDADFD6F7FFADDFE25896EE0198F96E159F2326208EB25B2D9FCC4B";
    attribute INIT_27 of inst : label is "EE320DFFF4CE67E7F9CB3FF0833E8FA6363ADE6F2BF6B36853E5FF35939FCFCE";
    attribute INIT_28 of inst : label is "FF17CA47787FA5557A87FA87F3F483343D98E0AD8000594E0AD80058E0ADD9CF";
    attribute INIT_29 of inst : label is "02FB869AFD1B26223A864BE8ECFD53027FF6DA12D3E5774457E394E001FACFBE";
    attribute INIT_2A of inst : label is "E7134942EEBBD37FAC9BCBB5EA75BFDF5FE96E23645FF44A7EBDBF02C4B12C08";
    attribute INIT_2B of inst : label is "37A9F70556BFE793D538F370ADFFC793AECEB91E4F8758BFA85AEB14AEC65012";
    attribute INIT_2C of inst : label is "4428EEFED4AC14A8100890894219FE11B47FCB37B5716A5B2FFF09FDDC748483";
    attribute INIT_2D of inst : label is "59B3FFF37FF9AE7FC100100000336FA40000020022DDBE9108080080000336FA";
    attribute INIT_2E of inst : label is "0003B968A1FFD8340B6E6FDFF258C86BF7F921AFDFF24B73C6DCD3FF67E9FBF7";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "4480009A49A410200281619494F40900200DBCC05E5423E525090A060AA22062";
    attribute INIT_01 of inst : label is "6641DE400E1601B04661700148800A0412806016058200142021080830909522";
    attribute INIT_02 of inst : label is "924DA1C4C2642999B24A46DA9890001BB59E6663B0002E6B0100200E6C2E072E";
    attribute INIT_03 of inst : label is "DA0559741016FF02050A05E33808A28005799484522B02089B9180F03C029265";
    attribute INIT_04 of inst : label is "FC58100B77EFF4FCDE1C1FF81FF818B65B2D16000015E6624C11818025AEEA0D";
    attribute INIT_05 of inst : label is "0E1285818008A1008114800EB620565F411D8025B2307C87F69E4018C006EFDF";
    attribute INIT_06 of inst : label is "080D8A70F114C4242881B14F914E42C3600ED29CC01025854480032C060013D0";
    attribute INIT_07 of inst : label is "68D7041F0D01800000000000800034EF514BA00084D03B91C00614885050C027";
    attribute INIT_08 of inst : label is "03CACB11CA28921C184571A6CFBA9B3200D3332517363B80C20DA0034C41303C";
    attribute INIT_09 of inst : label is "64592B2A00C6013C00C6E1045055FF0159801B846C88C0808DEEE47D9846C8BE";
    attribute INIT_0A of inst : label is "C4F8296B0011B8626213DD339802DB1610706047C600D639AC1557BF87294531";
    attribute INIT_0B of inst : label is "C7A180402C8B01C01F86C221C5F6ED8FE4605900BD08AEA01BC37052F20400E4";
    attribute INIT_0C of inst : label is "99749126C1015C649106C8A63B00FAECA8DDD6EC7C10012FD000A1EFC6400220";
    attribute INIT_0D of inst : label is "68268A62C8AD6546EEB763E138097E807EFFF8837AEF76770DE8919F65DD37BA";
    attribute INIT_0E of inst : label is "303252994612C140A6300883EC439AEDC8E1DF94F76FE1ECA9D7135BB7C937DB";
    attribute INIT_0F of inst : label is "000000C887000000CC21202248A588060000010331A0888818137BC061A0C001";
    attribute INIT_10 of inst : label is "240E00642400000000000000000B2810000005AA1056800D012C5A12502CA040";
    attribute INIT_11 of inst : label is "BA4400200AA0061601900034150300340804400CC0BC8000099200BCD2C05600";
    attribute INIT_12 of inst : label is "3330066400040000400940B1A4A068C04068308480B0B200AA00000B09A00AA0";
    attribute INIT_13 of inst : label is "54150541505415054150547FCFB1FFFFE2082AAAAA808A00005564AAABFFF333";
    attribute INIT_14 of inst : label is "100014A190468119046411505415054150541505415054150541505415054150";
    attribute INIT_15 of inst : label is "0000018A24202E842007C40802EA2408055543A481C5A110619081A2904054A9";
    attribute INIT_16 of inst : label is "0D48000C580018009050094540CB4D20C8033B6560000404CC07CC418309B481";
    attribute INIT_17 of inst : label is "2365A210243489428C0504009009428D00840080693EE0640CEDC01000008080";
    attribute INIT_18 of inst : label is "0A431000012B0003C4C8000DBD0B886AF802EA4100000D844020184077D2E874";
    attribute INIT_19 of inst : label is "0134E03E000F228034152589499600C00D06820034C884900222548000005000";
    attribute INIT_1A of inst : label is "6416841CDDDDCDDC406A411311244CCCCCD4B886B082C1166809030C18299034";
    attribute INIT_1B of inst : label is "991C21F9FBCC51C843DF3EC832E780555286B422AC2AAAAA83B11380FC19914B";
    attribute INIT_1C of inst : label is "283D1B1D0F56EB1987AB63C0F56C661E8D8F03D1B140F5643FDFBFDFE7BD5F5E";
    attribute INIT_1D of inst : label is "80102F56C56C18301E8DC09987AB23981E8C8D0F5646C87AB22643D1B1E87AB2";
    attribute INIT_1E of inst : label is "1003D1A00844400807B362801E8D00422200403D9B1E8D00422200403D9B1088";
    attribute INIT_1F of inst : label is "44400807B36289044400F4680211100201EED8C111003D1A00844400807B3631";
    attribute INIT_20 of inst : label is "8D00422200403D1B1888889044400F4680211100201EAD8A2224111003D1A008";
    attribute INIT_21 of inst : label is "90802662069A6D36C33468A82555E542B1555E5D7480F56EB19111112088801E";
    attribute INIT_22 of inst : label is "761821C30E3B1C76333DCB016CF4051EF81C5ACB3B984180551DB2040043675E";
    attribute INIT_23 of inst : label is "A4624460455480505804C10DA524166262E8240004400018CD920781C14C18F2";
    attribute INIT_24 of inst : label is "0420B30C16C821058A20B641082CD305B6084162082D90010A4010A4290A4290";
    attribute INIT_25 of inst : label is "0090821F600982184A483A00199B000382EE1195505A866104200084162082D9";
    attribute INIT_26 of inst : label is "0022633815A36000240000100010A59009FE00C2608692900B336824C2007052";
    attribute INIT_27 of inst : label is "1200A200001F884805104008D442700A56506824400B012AC40A81D047019191";
    attribute INIT_28 of inst : label is "00880195B4064262E5426540200234DCC059002D000004D002D00005002D1108";
    attribute INIT_29 of inst : label is "92C018007294900CCC5D16078800EB548008A0A408D1BA8888640D00000D0088";
    attribute INIT_2A of inst : label is "A024C4A4CBD15220C04D04D93CF80007E000A352DE1007A48000201480214970";
    attribute INIT_2B of inst : label is "C01202C9CE40C0430E3309637101984B004930612C0906D03266E8D1B09C52CC";
    attribute INIT_2C of inst : label is "B39001608A4B4BF1C9734BF32B25002427800221DFF27E6FB80040016B5A220C";
    attribute INIT_2D of inst : label is "A2E400003FE25C80010100000004905B400002020012006CA408080000000905";
    attribute INIT_2E of inst : label is "000014E63C004C98CE0508600B06065218002D486000A69D9DC1CA0005FF0205";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "DC3F098E51C81087D10D1FFBF10C4639280AB6801017A145B80D2E9307B31F13";
    attribute INIT_01 of inst : label is "4359CA962CA3BAF614B67E40B9F0100418009B96066E12143B32084803808560";
    attribute INIT_02 of inst : label is "388D0C95624D29AD94D286991CA5809B24DC545224BC789258C7184AA9815D2E";
    attribute INIT_03 of inst : label is "FA057F57D08106FA02763142B987B0029B689C6C00FB0086C59D2CA52944A0E9";
    attribute INIT_04 of inst : label is "879C1040BAB504284B9F2D52155AD8E4F279BD40A06DA2504FD92928200EEB0D";
    attribute INIT_05 of inst : label is "0D560800507068419C301F120618A9A0050FF080300E2C41D55A303FF0417562";
    attribute INIT_06 of inst : label is "7E0BC042D00094540A917809B8080AD07209E010C48624A1454BC29255E0F22E";
    attribute INIT_07 of inst : label is "E0104CBA1D1CDB6DB6DB6DB610000D6340C7A385592DBFB5C2E416A94938B80A";
    attribute INIT_08 of inst : label is "F0C2AA084608902E2C5145466A3B1B982C181109A11008F025975F86CE204174";
    attribute INIT_09 of inst : label is "3E630101E0EA0131E0B68D5B1F0D5FE015E003AB6A56CE196DEE8B7D1AB688AE";
    attribute INIT_0A of inst : label is "027F2A2831028162721211A9A47248100838301007F19C033A1555BDB7780455";
    attribute INIT_0B of inst : label is "A41CE27C27CC7178001680E1E0FECFCBA87C011CBD83BEBB12E25E50504800A4";
    attribute INIT_0C of inst : label is "964103E06A29733103C0608B21FFFB7E02BFD5FC48FB80E549E0E1555D782880";
    attribute INIT_0D of inst : label is "58C408B27CB1F015FEAFE245D4062A4F1E88F4C7EBE954450B4CC75759142568";
    attribute INIT_0E of inst : label is "99996ABD237C7EB2B5A1C383FC005E828A43DBBC556BC0840A52091374D62552";
    attribute INIT_0F of inst : label is "000001DF63000000417868281181984E00000001059B33301609C3CD44609E05";
    attribute INIT_10 of inst : label is "ED19811CD4F800000000000000052588000003A8209280A775290EEA5E149620";
    attribute INIT_11 of inst : label is "4A02842BAA5F01945FC900724D00C08C098C00E55F508D680358C0AB868BD405";
    attribute INIT_12 of inst : label is "3C380878000C001B40F2241049121220201000DB3F76B9225A0000076B9224A0";
    attribute INIT_13 of inst : label is "9A1589A1589A1589A1589A487005FFFFF575FDD555F7DD77772201DDDC889C3C";
    attribute INIT_14 of inst : label is "CC4A9922A00A001900A801589A1589A1589A1589A1589A1589A1589A1589A158";
    attribute INIT_15 of inst : label is "F870001D7B9C0EE39C6CA3E7C20E23E7C196652241E0A8CC090E713B0F3C18C8";
    attribute INIT_16 of inst : label is "25C9F834183E0602B7B06A8340F7D2302F87B796A005565457C099F600899DED";
    attribute INIT_17 of inst : label is "326461981D23A8860D0B3C007028860C000000001D2C2060C8B2CF8000008800";
    attribute INIT_18 of inst : label is "480EA3FF8118DF0089FDF079FD038F6AFF824BC03F0549BC4C3E1D5AD77CC465";
    attribute INIT_19 of inst : label is "400C6B9C0014238032D31FF25824A038220228F82BBD1964C5608B2CF810A3A1";
    attribute INIT_1A of inst : label is "1590B106DDDCDDDC404DEF8D9F770F0F0F122902291FAEC5BBDDE08B163FC972";
    attribute INIT_1B of inst : label is "4B2D39B1F304D8DE737F326C08486C4102A4850ACFFFFFFFC2A01421031E9445";
    attribute INIT_1C of inst : label is "E8018DF10073E8F98039BFF00637F800C6FC001CDF900637903510354AEB3F95";
    attribute INIT_1D of inst : label is "3A9820637F1224B600C69E878039BFE000C6FF0073FF08031FE1C01CFFF8031B";
    attribute INIT_1E of inst : label is "67524D7D4B199D4C1031BF3A926BEA58CCEA6081CDF26BEA58CCEA6081CDF633";
    attribute INIT_1F of inst : label is "199D4C0031BE320199D4935F52C66753040E6F80667524D7D4B199D4C0039BE6";
    attribute INIT_20 of inst : label is "6BEA58CCEA60014DF3232320199D4935F52C6675304086F8C8C80667524D7D4B";
    attribute INIT_21 of inst : label is "83037333F12C96596F3461FFFF01E10033F01F9933E004368F86464640333A92";
    attribute INIT_22 of inst : label is "4B2EF877CBA5874B1A2929C164FF851DFE1F4CFA2D120DF87D1BB06FC00887BF";
    attribute INIT_23 of inst : label is "A4CCAF810554EABBE039FFB62248573374B2907E02603C0E78D066F9779F2E4B";
    attribute INIT_24 of inst : label is "C521D8C91FEE290EC648FFF14876A047FB8A43B5823FDC29004010A4290A4290";
    attribute INIT_25 of inst : label is "0097E0155073FF6F4490AC8D9CDEBF2AE3FFBE1550AEEF742C81B8A43B5023FD";
    attribute INIT_26 of inst : label is "5C7BEB3F3FEBFC1480F82903E290A576295501BCFFDB91242BB9B224BFBF7802";
    attribute INIT_27 of inst : label is "0EBAA5DE051EC981F87C0C00760C5FF75B539031FC14818380CFF9F596995958";
    attribute INIT_28 of inst : label is "8F8C237BFC7F437B7484F485B3C2A37DFA9C9025000029C902D000289125104A";
    attribute INIT_29 of inst : label is "9D07BCDFDA8B242EE6165049B5E031741F0B6A8492E5FECDDFF25C9000020220";
    attribute INIT_2A of inst : label is "8F77F92C12CA45C02002022FB4EFAF38B0080A6FAA17842EE0A1AF1485214882";
    attribute INIT_2B of inst : label is "77BB828DF8F86E989B1BD3195DC0DE98851B1B7A62144E7F1A368285A1F640B6";
    attribute INIT_2C of inst : label is "508017CB8224C4DE465E46DE0CBE0134D4B8228EEA8A1425BF8340E1FD2CAC8B";
    attribute INIT_2D of inst : label is "EE00FE0AC00F409FC1100000000BE5D500000220003FD654600880000000FF59";
    attribute INIT_2E of inst : label is "000015289D7002FACFEFC1FF005FCE707F8109C1FE03EFBFD611D2F0920DFA0B";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "4C018BEC89CE88826F6A96DB253C0EB42C4A65231EF0525C2644E8D0E4E21041";
    attribute INIT_01 of inst : label is "514CC8C12A3356E6D1BBD140D335134610D0B2B30AC9151E2979A454311AC488";
    attribute INIT_02 of inst : label is "52EF2CD456821A1AC308602F3A104263614FE6EF5002769B07A13C2847870226";
    attribute INIT_03 of inst : label is "90D30BE42888030502689059DC88A8D3BC4E8271183D804A3C4F82D0B4201EA3";
    attribute INIT_04 of inst : label is "802A1522E221170A486CB912800A2BE3F0F8FC502AF13A28486484844C0851DB";
    attribute INIT_05 of inst : label is "2B489FE9150DB054D9460889E424F555090EC84F3E2101A27A52C99B4805C440";
    attribute INIT_06 of inst : label is "C906500469A025A60622CA80CA80101848978503E03EF141635021F73311C1B1";
    attribute INIT_07 of inst : label is "E003662F5C02DB6DB6DB6DB611040C6100C680416DB7A72660130E622A2844A8";
    attribute INIT_08 of inst : label is "08D231AC5242E70D0A300CE74FDD11EC02AB4B6AB4371990B7F278448351445E";
    attribute INIT_09 of inst : label is "7440FFFE102A019011F5762F4B5281131391434F543E776FE7E57F2AEDF55141";
    attribute INIT_0A of inst : label is "B460A3A3E89B3DC9FB010910384B638754342813C514F341E412395147C11548";
    attribute INIT_0B of inst : label is "4421CDC20E8809E63FE362D0303F532F35224092DE4B5F4480D0174343D02468";
    attribute INIT_0C of inst : label is "8E791624FA0128791604F2A893F77C71FF3BEDF3F1BF41E26A11613163440888";
    attribute INIT_0D of inst : label is "58D32A88E8918FF9DF6F9F8DDA0F13508F646880B457ABFD130881A2BBF44670";
    attribute INIT_0E of inst : label is "1B994AE573B46E96D4A026C1046034E28C61EDE0DA9DAC862027C5036E4E9803";
    attribute INIT_0F of inst : label is "000003CA220000006260701810802107000000C185400004033193B549548105";
    attribute INIT_10 of inst : label is "810500559784000000000000000300A0000001C40006A0C7A531CF4A600C0280";
    attribute INIT_11 of inst : label is "1AA8D60D2CC88503010500314742C4A883A11465F01166650EF2CAD7955F0B4F";
    attribute INIT_12 of inst : label is "C0380F8000097A2F50001410000A03B328519099401220A40A000001218A40A6";
    attribute INIT_13 of inst : label is "09114CD00489114CD114CD480004000010AA082AA88A80282828200A0A0A203F";
    attribute INIT_14 of inst : label is "FF715FD7305001620500122401114CD22401114CD22401114CD22401114CD204";
    attribute INIT_15 of inst : label is "0522AA8087FE48C7FE6BC7FFE5E1E7FFE6186127E60645FF545FF93B9FFF610D";
    attribute INIT_16 of inst : label is "212084570C11140824142001D0259B14A85CACD4608542429C25AD484280893D";
    attribute INIT_17 of inst : label is "76D56560496914038401B00120140384004000485180843469FAE80000000004";
    attribute INIT_18 of inst : label is "1305AD60C5539082D3490859BC874D29C8401D0510851B7104610A225DDF4E3E";
    attribute INIT_19 of inst : label is "4086720C0004588018518580894E50B16B2479841979EDF5FE2AE93D805025E9";
    attribute INIT_1A of inst : label is "24668D94DDCDDDDC5A183EBDF294700FF01C784630A17EE6B4A512848E210531";
    attribute INIT_1B of inst : label is "9286296C0F9DA47C52E0FBD21298B73ED48B3480F47FFFFFE4CC941105C9514F";
    attribute INIT_1C of inst : label is "2A00D5118035631E401AA308025461006A8C200D511802546AE5EAA5CCCDAAB3";
    attribute INIT_1D of inst : label is "056C2025C70183B1004BF180401AE201004B8F802547FC01AA3FE00D518C012A";
    attribute INIT_1E of inst : label is "00AC41E2B20002B60012E205620F15900015B080D7120F15900015B080971400";
    attribute INIT_1F of inst : label is "0002B6001AE20010002B1078AC8000AD8406B884000AC41E2B20002B6101AE20";
    attribute INIT_20 of inst : label is "0F15900015B08017100000010002B1078AC8000AD8002B8800004000AC41E2B2";
    attribute INIT_21 of inst : label is "51D15555092DB6496FB46005C001E14030001E1EF068005E3100000002000562";
    attribute INIT_22 of inst : label is "9A94F4A7A54D4A9AAA2E6EA443B04934691A0EE6AD97454468489A2A2100CD1A";
    attribute INIT_23 of inst : label is "B4514110055791501C2D76DE8F7BD11115FE00E1324512347CDA33C4A7DE945B";
    attribute INIT_24 of inst : label is "24A97A000DB8254BD0006D492A5E10036A0952F0801B5285214850B52D0B52D0";
    attribute INIT_25 of inst : label is "9680028A285AEDBD1EF7BFA40445F097D19D045558BE4B5500A080952F4101B5";
    attribute INIT_26 of inst : label is "6A5ED3EBFB7AF210B444215112D4B40828A28736BB6F07BFE888FE8275F0CE5A";
    attribute INIT_27 of inst : label is "04D2D4F10449E0E08659060A4505F8126367D8916A1EC42070678526FDF45455";
    attribute INIT_28 of inst : label is "E0461ED2CFD9511195BC95BEDE288F776410527D000040C527D00040535D767B";
    attribute INIT_29 of inst : label is "15252FEDBC3FBFE2229FC4C93792184608827A249225665444414C50010B3673";
    attribute INIT_2A of inst : label is "B294C044A760E090B06A14AAA64E80AC282288DC821041829081208280A82978";
    attribute INIT_2B of inst : label is "694A48ACA1443FFAA3C8FE5BDF2047F2CE294F1FCB3885706BD55AF5585FC0D6";
    attribute INIT_2C of inst : label is "F4385F8F90E71E9D1C1D1C9C4DF410F6D184084B88838524D8474012E76FBFEF";
    attribute INIT_2D of inst : label is "FAB0410A400ACE0800000000002FF78F0000000000BFDF3D0C0000000002BE78";
    attribute INIT_2E of inst : label is "0002450ED90803B4FAD468F0896F7CCA3C478328F10FEDF25E049A0880060502";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "282950400C2A188AF2420C025CD0812408E0840B9A010D5D780CF01A0AA44446";
    attribute INIT_01 of inst : label is "783888C4303826110304C8572F5C9D060D4303E3040F1F060D608C7C15484008";
    attribute INIT_02 of inst : label is "512A10A4A4C2101102084C8A781114E4E949808FA06962A209488408750A0874";
    attribute INIT_03 of inst : label is "055A8062828028D0AC3992009082714610090450085180142009080000129125";
    attribute INIT_04 of inst : label is "810D4CA00205152848C93152355293E5F3F9FD4A49402409010901014AB01452";
    attribute INIT_05 of inst : label is "28805022221B173340400C2A4E52A5AA130251525C482C0DBABA21D885200402";
    attribute INIT_06 of inst : label is "8851800C098021B6042230014001004D6802200100E152004242946002A48044";
    attribute INIT_07 of inst : label is "4987503AB811C924924924922140B5EC81CE020C9449338420803642281020E0";
    attribute INIT_08 of inst : label is "A1DAE3389A7FC6DED42965956A9F5B1420C3736C373653054A04852145634831";
    attribute INIT_09 of inst : label is "8C9B5554C512B80D4586C298A80DC04392056260754109901017608E8E0F4561";
    attribute INIT_0A of inst : label is "A5443333200BB4FAEA994998B5524306DB7B5358124CA7C14F0AB9E9E041F559";
    attribute INIT_0B of inst : label is "EDF204A8F1936313751147301F395B622C106480C20CD1406DEDA8424240048A";
    attribute INIT_0C of inst : label is "16441F2F00323C841F0F0EAABC20845155AA2D53404515001145013503114079";
    attribute INIT_0D of inst : label is "7AC0EAAB191C8AAD516A9A0200A9008A5108A901A64976450F79073259153DEA";
    attribute INIT_0E of inst : label is "060614114042013CA72114002C1428C2AE6228209B0AA3DC0377611FE41E055E";
    attribute INIT_0F of inst : label is "00000210C4000000091908004127B9C0800001E0202000015C6073A81C275438";
    attribute INIT_10 of inst : label is "0260862724500000000000000008A8580000042000BC87C04A37C0946822A160";
    attribute INIT_11 of inst : label is "B264B07A4D34281214D4800538944780791132449AA4010C58B020B483F21A19";
    attribute INIT_12 of inst : label is "FFC00000000021524ABB52A5BDA96D10E28864C60AA01A92A200000A00292B20";
    attribute INIT_13 of inst : label is "09916CD916CDA2601A2601C8000600001D57D5DDDFF75D5DF75DE7D77DD7603F";
    attribute INIT_14 of inst : label is "019DE01B306001B306CC180601916CDB36CDA260180601916CDB36CDA0609806";
    attribute INIT_15 of inst : label is "A9B4CD1F500088C800C288001B1618001FEF9ED81A5FFE01F7600233A000FFF2";
    attribute INIT_16 of inst : label is "7524D186849C40104140030625CBE1334D3A33271229868626928A7114519489";
    attribute INIT_17 of inst : label is "36400470305621C001060800C021C00100940092882CB30060B4B50080080001";
    attribute INIT_18 of inst : label is "19261AD494690A2853C8A2AB02A9AA110D174E281A29192005B452327576CB66";
    attribute INIT_19 of inst : label is "213A89A0000902000606A87100382510C01C3A5146591691533F26F1509502E6";
    attribute INIT_1A of inst : label is "76C2944A9899999802CDF34BEE767FF0000EF41C7C5F1355779DC40A0380D485";
    attribute INIT_1B of inst : label is "4902495C0BF8803092A0BD814857700DBD981580C2D7FFFF911DC7D600059C4B";
    attribute INIT_1C of inst : label is "A8E9F9D13A7E49D81D3F3B03A6E76074DCEC0E9B9DE3A7E71595159570F1CCDA";
    attribute INIT_1D of inst : label is "C001AA7E7500004E74DCCC801D3F3A0074DCED3A6E7609D373A04E9B9D89D3F3";
    attribute INIT_1E of inst : label is "F801BE0005FFE000C5373BC00DF0002FFF000629B9DDF0002FFF0006A9B9DBFF";
    attribute INIT_1F of inst : label is "FFE000C5373BFFCFFE006F80017FF800314FCEF3FF801BE0005FFE000D53F3BF";
    attribute INIT_20 of inst : label is "F0002FFF00062979DFFFFFFCFFE006F80017FF800354BCEFFFFF3FF801BE0005";
    attribute INIT_21 of inst : label is "01117777A04104004B4B9FFA3FFE3EBFCFFFE5E00F93A5E49D7FFFFFF9FFC00D";
    attribute INIT_22 of inst : label is "434CFA67D321A6435A2909C571220E64083F8162211405E0FE68502F0ACDC902";
    attribute INIT_23 of inst : label is "A0550410055504144144B0A08481137372808A943841104C081032E2679F4C42";
    attribute INIT_24 of inst : label is "850382411FEC281C1008FF6940E09047FB4A0704023FD900001004A0280A1284";
    attribute INIT_25 of inst : label is "8002A02082896141090220020DDD4A42E3FF105552C2CB78310294A0704023FF";
    attribute INIT_26 of inst : label is "54B15D80C7D3F8A0125140C9400400A202002E425850424089BB800A014A7800";
    attribute INIT_27 of inst : label is "3BA4C3485800C0A4D21C04AC45265D041C16005070B00AB2526353F50C6A9A9B";
    attribute INIT_28 of inst : label is "2ACD4495C1144331C5504511254982F1744D4D0100004414D090004548091140";
    attribute INIT_29 of inst : label is "0288955402124086EE5001450A427C440C28948210FDEEDDDD35214800501820";
    attribute INIT_2A of inst : label is "BE7738801C18042513A1184D46DE2A10B295E66C0355140EC5323A9400080080";
    attribute INIT_2B of inst : label is "EF3B0AAEA961F3416FF9E8257E8BCF494C297C3D253085EAD3A550A157F0DAAE";
    attribute INIT_2C of inst : label is "929039400A420A1A0A9A0A1A28F866B724B179440A8A9424152A7AA7FD5C324A";
    attribute INIT_2D of inst : label is "C2005453C003424A80000080089890490200200000624124A40000040045C904";
    attribute INIT_2E of inst : label is "0000552B1042BC576038C0FA151533803E0ECA00F85D825F11580AA29055D055";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "582752A94ABC51971A028480561405A09AC9FE933440B6A072CCB9B7D7B64545";
    attribute INIT_01 of inst : label is "600DAACEBC700EA980204AE429143A2C508826AE289A363C7B0D18D893910801";
    attribute INIT_02 of inst : label is "150952A4E656B511924A5E3A5A93A46A2C58090A4225AB84355A053A450125FF";
    attribute INIT_03 of inst : label is "48DEC1C254E3C4CA900870A1719CF08914784210111F1034085B1DA368D29525";
    attribute INIT_04 of inst : label is "7A7D200D7F4AECD5FD793FAB7FFBDAF5FAFD7F6C8051E12020FB1B1A691636D6";
    attribute INIT_05 of inst : label is "A8C0BD8401E7258040445D63AA3A0500D526D51D4C0AFCD7A23455F294CAFE9D";
    attribute INIT_06 of inst : label is "1A908939E2124B2C84881127012707EBE022A24E4888D411CA464404A1888192";
    attribute INIT_07 of inst : label is "4DB7D05A4874B6DB6DB6DB6CF40AB5EF1B5FC6AA024977D4C8A2B648A8B06AB4";
    attribute INIT_08 of inst : label is "95DAEB3ADA62B6DEDD656D9D5A73FB4434C36A6C36A67719410414A85B6BF9B2";
    attribute INIT_09 of inst : label is "AECDD5D4A95A1207298C51386A30802B39295730D4A12856121D709AB90D7BC1";
    attribute INIT_0A of inst : label is "954D2B2B6443335150C7BC7733F24B56DB7B753FE02EBAFD772228D0E0E34BB4";
    attribute INIT_0B of inst : label is "8888BFE575D9D5481567D6E64469E29BE1755E25B3ABB9E86DEDBA5A5AC0151A";
    attribute INIT_0C of inst : label is "B0C6D3704DABB126D3504977010243D554323996D7412514832961CAA18A7382";
    attribute INIT_0D of inst : label is "5B1497715DD6AAA191CCB6BA2128A4197199CD89B25822C76BDD9F92C31DAF7B";
    attribute INIT_0E of inst : label is "50501109DA1B4B30E5135E0825DB81DFDDE63C31AA193AB4E33F57666418A7C7";
    attribute INIT_0F of inst : label is "FFFFFC2008FFFFFF100207C1041FFFF07FFFFFFC4200000255E54561028032A0";
    attribute INIT_10 of inst : label is "024210A4254BFFFFFFFFFFFFFFF04207FFFFF8114E0016D408B5A8116BC1081F";
    attribute INIT_11 of inst : label is "403199684C954A0212207F8800250450C56001F4B902108895B4001DE1520A09";
    attribute INIT_12 of inst : label is "00000000000D5040C48081CE0040824014A10AA24908440840FFFFF084408400";
    attribute INIT_13 of inst : label is "CC220000008800000330CC480001FFFFE22A00A0A0A80A8A2820A00820A2BFC0";
    attribute INIT_14 of inst : label is "FE6600033000003300CC0330CC22000000000000000000110CC330CC310CC310";
    attribute INIT_15 of inst : label is "9E00F1AAAFFF08D7FF7737FFF4C997FFF7FFF7E7E5A7F9FE089FFCC45FFF0005";
    attribute INIT_16 of inst : label is "6D83CA87587A886040838438094B840A4CA12926004FC1C1A652AA602500424B";
    attribute INIT_17 of inst : label is "B440826F8200403853F043FE0FC03853FF0FFF04A6108805E2F4948080800002";
    attribute INIT_18 of inst : label is "061D1853A550A949CB0A94A183B56A772CA69A11794F11201E32D9BF08800887";
    attribute INIT_19 of inst : label is "1E410001FFE0845FC10840042201094114016D4A42DFC04B212052EB483958A3";
    attribute INIT_1A of inst : label is "9172924ECDDDDDDC428EE9239EF680000012C2284A2708347BBDA50A42C22008";
    attribute INIT_1B of inst : label is "384362868703BA3AC528701C79F8837A71899336DA280000155DAC43FCD85CA9";
    attribute INIT_1C of inst : label is "697D41B15F4059BFAFA837F5F506FEBE80DFD7D41BF5F406BF0BBF4BC0FE0F1C";
    attribute INIT_1D of inst : label is "ED728F506C7FBF7EBE80AAFFAFA037FEBE80DD5F506DFAFA037F97D41B82FA03";
    attribute INIT_1E of inst : label is "FDAE7FE6BB3FF6B957A037ED73FF35D9FFB5CABD41B3FF35D9FFB5CABD41B67F";
    attribute INIT_1F of inst : label is "3FF6B957A837FFB3FF6B9FF9AECFFDAE51EA0DECFFDAE7FE6BB3FF6B957A036F";
    attribute INIT_20 of inst : label is "FF35D9FFB5CA3D81B7FFFFFB3FF6B9FF9AECFFDAE55EC0DFFFFECFFDAE7FE6BB";
    attribute INIT_21 of inst : label is "1797777796936934923B7FEE7D7453B687D740FFF7C5F6059B8FFFFFF67FED73";
    attribute INIT_22 of inst : label is "E35DFAEFD771AEE37AAB8BD56B62AC6E1ABF3162B15C5DEAFCFC72EF531A9BC6";
    attribute INIT_23 of inst : label is "00FFFAB15003EEFBE273F58DDDA6137372CC3552B4C1755D8B12EBEAEFBF5D62";
    attribute INIT_24 of inst : label is "C106A3ED9FEF08351D6CFF7841A8EB67FB820D47DB3FDDA86A0A840000401000";
    attribute INIT_25 of inst : label is "9417E29544E7EB1ABB4C330DCDDF2963E3F7EAC00412DB7C2F854C20D47DB3FD";
    attribute INIT_26 of inst : label is "C4FE7DD20FE3F93065CA60172284A176295448D9FAC6EED309BBCC279A297850";
    attribute INIT_27 of inst : label is "AA84D12A9C01C3C3CC101D39C61D7C80808920B8412105EA21FF4BFC4F0B3B1B";
    attribute INIT_28 of inst : label is "598C5DB5E2327331A76327226D0988F3702204587FFF82204587FF8200702BD4";
    attribute INIT_29 of inst : label is "BF9E7F457776D306EE5984E5D96A7AC43D44A68049FDEEDDDC880207FE94177D";
    attribute INIT_2A of inst : label is "4EF60211000408094054254F7C1C395744EA34F8660CB75EE9AB019425094152";
    attribute INIT_2B of inst : label is "F77BAAACA569E826273985CD7A93CC2E5C29BA30B97087E9224568D153D8368E";
    attribute INIT_2C of inst : label is "9290231DCA664E5E4EDC4C5C2EFEAAB5476A4035FD766AFEF488C08FFD5E2928";
    attribute INIT_2D of inst : label is "E321F29F3C035C3E500000808015AEB9020200000046BAE4A480000404015AEB";
    attribute INIT_2E of inst : label is "000154E670D4D39F74980BF95B808282FEA8AA0BFA90B69E99D00994FF88CA95";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "BE3FD9447664808F9918364B341A07904FCCF47F0153DF44199509733DE26773";
    attribute INIT_01 of inst : label is "4B938B37FFB1986111925FFD99257A502E959F22127E04001FB928186FB28480";
    attribute INIT_02 of inst : label is "018018333C0631EE5D75BC8918EDFDB1009A66623DBF9E33D1FBDC03AD87DA2C";
    attribute INIT_03 of inst : label is "726FFC13EFEE80FDF6F871411B8F1E94DC68897010E108F20411EF5DFF7CE198";
    attribute INIT_04 of inst : label is "878FF015FAB500280B8FCD54F554F0A05028149F9271A230878EEFEFDC44BE67";
    attribute INIT_05 of inst : label is "F148E903B1F1052118443FE4A03F5655C40B7F652A3F837D766BBEB17FDBF562";
    attribute INIT_06 of inst : label is "07F276CCA86DA08206A44E999E991248208B3D30A09034402353FC921FFEC6AF";
    attribute INIT_07 of inst : label is "32091105049E92492492492511A7C252242513FC4B649E94A0FDF66A0A69BFA0";
    attribute INIT_08 of inst : label is "FCA514C6218889CBC7B082044D121B0C4F1C9991C99999FF6DB25FEDC73F0A08";
    attribute INIT_09 of inst : label is "9C432B2BFF6A9911FF32C10BDB1DC3FF00FFC0233E068C18681FC35FC233E161";
    attribute INIT_0A of inst : label is "106F8C8C0214C55151C10810C4392C19CF2F1FC839E27A04F7977C64792CC31C";
    attribute INIT_0B of inst : label is "841E603FF3887F3D8A93FE304C71D4CFA43FC49FD3F8D9FCE4BC8F191800BE8E";
    attribute INIT_0C of inst : label is "186C71F138E1739C71C1386384A84364AC843C266B447CA541FFC015047FE590";
    attribute INIT_0D of inst : label is "9405863938B1256421E1335A0BE42A0FD08898A3E2CD76699A50A11661A6694C";
    attribute INIT_0E of inst : label is "090B1A242124259610E1F2216E78044584321A765F4E7E952475C0955AE02D64";
    attribute INIT_0F of inst : label is "000003DFF7000000EFFDF83EFBE0000F80000003BDF80007C320C16428C05FEC";
    attribute INIT_10 of inst : label is "89030931907C000000000000000FBDF8000007EEB1043E432514865A2E3EF7E0";
    attribute INIT_11 of inst : label is "008853E124CFFB1E1FDF8077FFFD841841A005C60FFDEF7BF6E0D0B607CB1E05";
    attribute INIT_12 of inst : label is "FFF80FFC000D7BCB06FF7E31FFBF7E610FB080810FF7BBF41000000F7BBF400C";
    attribute INIT_13 of inst : label is "0080200A220080200B32CCC80003FFFFEAA0AA00AA000A0A802A200A80A83FFF";
    attribute INIT_14 of inst : label is "FE80200B302000B302CC0B32CCB32CCB32CCB32CCB32CCA22008020082200822";
    attribute INIT_15 of inst : label is "F007018AAFFEB10FFE800FFFE8000FFFE8000FEFE80FFBFE803FFA003FFE8003";
    attribute INIT_16 of inst : label is "E403FF91087FEC6027FC7BC7FF25B60267EC8DB3F2FC424293FC033FFD800B24";
    attribute INIT_17 of inst : label is "2E20C1A87DFFBFC7AC0FBC01F03FC7AC00F000FFB4145021E0B64F8088000007";
    attribute INIT_18 of inst : label is "021DC97FFE359FFCC0C1FF9881810123BFFE43107FFC18B01C1FCA38A8226437";
    attribute INIT_19 of inst : label is "E1BEFFFE001F7BA03EF7BFFBDDFEFF600630087FC96489248D10D964F87F3129";
    attribute INIT_1A of inst : label is "198CBBF2202220220FC4248D82137FFFFFF2A3782B012580B084FD8BE687DFF7";
    attribute INIT_1B of inst : label is "07C620B483040E6041483047D6C86C38700C6840C78000003C4CF04D0F0E1B04";
    attribute INIT_1C of inst : label is "F7E84CF1FA1306FFFD019FFFA033FFF4067FFE84CF6FA133F575F535FF000FE0";
    attribute INIT_1D of inst : label is "EFFF8A133FFFFFFFF4263F807D019E01F40678FA133FF7D099FFBE80CF07D019";
    attribute INIT_1E of inst : label is "FDFF7FF7FFFFF7FFD5099FEFFBFFBFFFFFBFFE284CFBFFBFFFFFBFFE280CFFFF";
    attribute INIT_1F of inst : label is "FFF7FFC5099FFFFFFF7FDFFDFFFFFDFFF14267FFFFDFF7FF7FFFFF7FFD5019FF";
    attribute INIT_20 of inst : label is "FFBFFFFFBFFEA84CFFFFFFFFFFF7FDFFDFFFFFDFFF14267FFFFFFFFDFF7FF7FF";
    attribute INIT_21 of inst : label is "07871111F92DB6CB2E7FFFFF7FFEF7FFD7FFEDFFFFFFA1306FDFFFFFFFFFEFFB";
    attribute INIT_22 of inst : label is "19C43E21F10CE219D80860FE2073FD0C5FF3044004161C7FCC38F0E3FF3803B6";
    attribute INIT_23 of inst : label is "001100100001151457CC731606C8C5151832123FF0007FC42040E2FE2187C458";
    attribute INIT_24 of inst : label is "D00E5E582B278072F2C159340397860AC9A01CBCB0564E004000020080600802";
    attribute INIT_25 of inst : label is "4002A0200F98E62D0D918C8494449FCAF59100400F6F4714648CBA01CBC30564";
    attribute INIT_26 of inst : label is "0FB9B99962D8BFD1A1FFA307E80200220200FB26398B43646288B202649FCD00";
    attribute INIT_27 of inst : label is "E612449FF408C3CBFCCE1FF8025C5FFF7F79B1133FE588A005CBFF3098BE4E4F";
    attribute INIT_28 of inst : label is "0F87C6E2C8D92557908D90CC97FF8370FFDDFA2800007DDFA200007DFE005421";
    attribute INIT_29 of inst : label is "22B98D8CDA19646A230640506CFF18003FF65A0DB66C774447F7FDF801F63000";
    attribute INIT_2A of inst : label is "8213FDEEFFFBF7FF60260264F44DEFCEBFE8662C22B7FC027EEDEF4030040000";
    attribute INIT_2B of inst : label is "6109FC04C87F64B18B1A963118FED4B9C0091952E700046F8910664C1EC60017";
    attribute INIT_2C of inst : label is "C8C86C86A309615B63DB635B8139FE109C3FE013EA8014051FFB06FDCC2C8583";
    attribute INIT_2D of inst : label is "C9E1FFF9C0193C3FC00000880032430C0220000000C94D323000000440036430";
    attribute INIT_2E of inst : label is "0003E33A037FD26E6648C3BFF908D800EFFB8003BFF6CB724740A6FFF500FDF2";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC093C7700020300";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "F83FDBCC46E4000F9B18365B340C03B12FC4407D1043FE00398407F137C12721";
    attribute INIT_01 of inst : label is "49510A07D6131AC130B24FFD99283A141E859F44167C08043F39002007B08400";
    attribute INIT_02 of inst : label is "018118307A042106D14638933081FDC642166266103F9E1110F9D80209851E28";
    attribute INIT_03 of inst : label is "623CE443FF6E82FFF6C07001238F3E85DC00896010C200F204108FF1FC718180";
    attribute INIT_04 of inst : label is "0397F015C810040061938000E008E8804020101F90700230439F8F8FB454A634";
    attribute INIT_05 of inst : label is "D9C0F9021072052108043FEEA23F5255C4003F35020F807844E03F91BFDB9020";
    attribute INIT_06 of inst : label is "17F24002C400114506104800080002C84009B000C08040004343FC9231FEC0AF";
    attribute INIT_07 of inst : label is "00110005201E36DB6DB6DB6C30078043000583FC4B258688C4F1E66108303FA2";
    attribute INIT_08 of inst : label is "F88018844108918B8FD00004472036080E0800008001E65F25B2CFED8A3F0009";
    attribute INIT_09 of inst : label is "B82A2A2BFF3A0005FEB08113D1193CFD117EC3231A068408681983531031889E";
    attribute INIT_0A of inst : label is "004F88880030055151C21021043928118E2E3FC83BE74C469B044E86B828C304";
    attribute INIT_0B of inst : label is "029EE4FFD7057E7C0A81BE004C4180C4041FC00F03F8019CC0B81B1110013B80";
    attribute INIT_0C of inst : label is "882C70F178E043BC70C1786105AAC304A840320420407C8401FE6150013FE590";
    attribute INIT_0D of inst : label is "F00D8611702425420190210223E5200F80801042C084442C1630400420B058C0";
    attribute INIT_0E of inst : label is "191B1824632464921181E60048780C87084210740C4444002052C10CCA80683C";
    attribute INIT_0F of inst : label is "000000000000000000000000000000000000000000000007C741814400C01FEC";
    attribute INIT_10 of inst : label is "89030010907C000000000000000000000000000000103E062C040C580E000000";
    attribute INIT_11 of inst : label is "008853E160DFFB041E000000007D8498C9E001C50F00000BF6C1D0260C9B040D";
    attribute INIT_12 of inst : label is "FFF80FFC000D5BCB04E00000000002602FB010830F0000000000000000000000";
    attribute INIT_13 of inst : label is "000000000000000000000037FFF9FFFFE02AAAAA00000AA0002A82A000AA9FFF";
    attribute INIT_14 of inst : label is "FE001FE000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "F007FD8AAFFE39C7FE7FE7FFE7FFE7FFE7FFE7E7E7E7F9FE7F9FF9FF9FFE7FF9";
    attribute INIT_16 of inst : label is "E003FFB3007FEC20278000001F64B61227E48C9200FCC0C093F003207DC0092C";
    attribute INIT_17 of inst : label is "2900C1C00000000000000000000000000000000FB0104201C0920F8000000007";
    attribute INIT_18 of inst : label is "021DA17FFB1ABFFA00A3FF944101211227FE21007FFC04301F1FC45A20822415";
    attribute INIT_19 of inst : label is "00000000000000000000000000001F602600087FCB648B248C00CB2CF87F3123";
    attribute INIT_1A of inst : label is "1190BBC6020022200DA42C8C923300000010AB7A23012C91908CFD83E6060000";
    attribute INIT_1B of inst : label is "00C0109483001E082108300FD0980010508080024B8000003800704F00061804";
    attribute INIT_1C of inst : label is "E3C044FFF01108F078089E0F0113C1E022783C004F8F0013E060E060FFFFF000";
    attribute INIT_1D of inst : label is "FFFF80113FFFFFFFE0223FFFF8089FFFE0227FF0013C0F8009E07C004FFF8009";
    attribute INIT_1E of inst : label is "FFFFFFFFFFFFFFFFC0089FFFFFFFFFFFFFFFFE0004FFFFFFFFFFFFFE0004FFFF";
    attribute INIT_1F of inst : label is "FFFFFFD0089FFFFFFFFFFFFFFFFFFFFFF40027FFFFFFFFFFFFFFFFFFFC0009FF";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFE8044FFFFFFFFFFFFFFFFFFFFFFFFFF40027FFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "07871111F92DB6D92FFFFFFFFFFFFFFFF7FFFFFFFFFF00108FFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "49C41E20F124E249C80920FB2143F42817F30C400C121C7FCC7060E3FF380AA4";
    attribute INIT_23 of inst : label is "001100100003001507CC221682D8C1111412127FD0407FC460C0E27E2083C448";
    attribute INIT_24 of inst : label is "E00E48400966007242004B300392100259801C900012CF000000040100000000";
    attribute INIT_25 of inst : label is "0002A0000F98442D05B184848445BFDA719100400F26411C01803C01C900012C";
    attribute INIT_26 of inst : label is "0F99A99122489FF021FFE007F00000AA0000F966110B016C6088921065BFCE00";
    attribute INIT_27 of inst : label is "EE1605BFFC0043C3FCC21FF8421C4F800008B00303ED802001E97F30B09E4E4F";
    attribute INIT_28 of inst : label is "0F87C2C258C92111118C918D97F4833038000000000000000000000000004421";
    attribute INIT_29 of inst : label is "00B984889A096C622282404865FD18403FF24E00002466444780000001F61000";
    attribute INIT_2A of inst : label is "023300000000001F60260224C0258FCE1FE865242007F0067F8F8F0000000000";
    attribute INIT_2B of inst : label is "2119F604087F2CB18908963108FE44B988090B12E620042F993022440E421232";
    attribute INIT_2C of inst : label is "C4A865869299514B53CB534B4319FE30B03FE0132002003027FB04FCC4258D83";
    attribute INIT_2D of inst : label is "4921FFF90019243FC00000000036D34C0000000000DB0C312800000000032C30";
    attribute INIT_2E of inst : label is "0003B002107FD26A6448039FF908C800E7F980039FF2D932420050FF7505FFF2";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1D1C7600000300";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
