library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_PROG_ROM_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_PROG_ROM_2 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"CA",X"CA",X"10",X"E1",X"A5",X"43",X"30",X"0E",X"C5",X"42",X"90",X"0A",X"69",X"02",X"C9",X"1E",
		X"90",X"02",X"A9",X"FF",X"85",X"43",X"A6",X"CE",X"30",X"05",X"A0",X"4F",X"20",X"16",X"77",X"A9",
		X"00",X"85",X"22",X"85",X"41",X"60",X"86",X"0C",X"8A",X"4A",X"AA",X"94",X"42",X"84",X"10",X"C4",
		X"CE",X"B0",X"26",X"84",X"CE",X"A9",X"00",X"85",X"11",X"98",X"38",X"E9",X"03",X"90",X"04",X"E6",
		X"11",X"D0",X"F7",X"A5",X"11",X"49",X"FF",X"69",X"04",X"85",X"11",X"06",X"11",X"65",X"11",X"06",
		X"11",X"65",X"11",X"85",X"CC",X"A9",X"14",X"85",X"CB",X"A2",X"1B",X"E4",X"10",X"F0",X"1D",X"B5",
		X"41",X"95",X"44",X"B5",X"42",X"95",X"45",X"B5",X"43",X"95",X"46",X"B5",X"20",X"95",X"23",X"B5",
		X"21",X"95",X"24",X"B5",X"22",X"95",X"25",X"CA",X"CA",X"CA",X"D0",X"DF",X"A9",X"0B",X"95",X"44",
		X"A9",X"00",X"95",X"45",X"95",X"46",X"A9",X"F0",X"85",X"77",X"A6",X"0C",X"B5",X"64",X"99",X"25",
		X"00",X"B5",X"63",X"99",X"24",X"00",X"B5",X"62",X"99",X"23",X"00",X"4C",X"FF",X"6F",X"98",X"10",
		X"09",X"20",X"B6",X"70",X"20",X"AA",X"70",X"4C",X"B6",X"70",X"A8",X"8A",X"10",X"0E",X"20",X"B6",
		X"70",X"20",X"BC",X"70",X"49",X"80",X"49",X"FF",X"18",X"69",X"01",X"60",X"85",X"0D",X"98",X"C5",
		X"0D",X"90",X"0E",X"A4",X"0D",X"85",X"0D",X"98",X"20",X"D1",X"70",X"38",X"E9",X"40",X"4C",X"B6",
		X"70",X"20",X"EB",X"70",X"AA",X"BD",X"D9",X"70",X"60",X"00",X"02",X"05",X"07",X"0A",X"0C",X"0F",
		X"11",X"13",X"15",X"17",X"19",X"1A",X"1C",X"1D",X"1F",X"20",X"D5",X"A0",X"04",X"C5",X"0D",X"90",
		X"02",X"E5",X"0D",X"26",X"0C",X"0A",X"88",X"10",X"F4",X"A5",X"0C",X"29",X"1F",X"60",X"18",X"69",
		X"40",X"10",X"08",X"29",X"7F",X"20",X"0B",X"71",X"4C",X"B6",X"70",X"C9",X"41",X"90",X"04",X"49",
		X"7F",X"69",X"00",X"AA",X"BD",X"61",X"4B",X"60",X"A9",X"04",X"85",X"76",X"20",X"A2",X"4B",X"C6",
		X"76",X"D0",X"F9",X"A2",X"C9",X"A9",X"47",X"85",X"04",X"A9",X"02",X"85",X"03",X"A9",X"C1",X"20",
		X"D5",X"7C",X"A9",X"BE",X"85",X"09",X"A9",X"75",X"85",X"0A",X"A9",X"00",X"85",X"01",X"A9",X"70",
		X"A2",X"20",X"20",X"7F",X"71",X"4C",X"D6",X"79",X"A9",X"C5",X"A2",X"C9",X"20",X"D5",X"7C",X"A2",
		X"BE",X"A9",X"75",X"85",X"0A",X"86",X"09",X"D0",X"2E",X"AD",X"03",X"28",X"29",X"03",X"A2",X"10",
		X"86",X"01",X"0A",X"AA",X"BD",X"F1",X"71",X"85",X"0A",X"BD",X"F0",X"71",X"85",X"09",X"71",X"09",
		X"85",X"09",X"90",X"02",X"E6",X"0A",X"98",X"0A",X"A8",X"B9",X"D4",X"71",X"BE",X"D5",X"71",X"20",
		X"1F",X"7A",X"A9",X"70",X"20",X"EA",X"7A",X"A0",X"00",X"A2",X"00",X"A1",X"09",X"85",X"0C",X"4A",
		X"4A",X"20",X"B0",X"71",X"A1",X"09",X"2A",X"26",X"0C",X"2A",X"A5",X"0C",X"2A",X"0A",X"20",X"B6",
		X"71",X"A1",X"09",X"85",X"0C",X"20",X"B0",X"71",X"46",X"0C",X"90",X"DF",X"88",X"4C",X"55",X"7A",
		X"E6",X"09",X"D0",X"02",X"E6",X"0A",X"29",X"3E",X"D0",X"04",X"68",X"68",X"D0",X"EE",X"C9",X"0A",
		X"90",X"02",X"69",X"0D",X"AA",X"BD",X"F6",X"56",X"91",X"03",X"C8",X"BD",X"F7",X"56",X"91",X"03",
		X"C8",X"A2",X"00",X"60",X"68",X"B6",X"72",X"B6",X"0C",X"AA",X"0C",X"A2",X"0C",X"9A",X"0C",X"92",
		X"68",X"C6",X"6E",X"A7",X"56",X"42",X"5A",X"42",X"58",X"42",X"68",X"32",X"64",X"C6",X"6E",X"D2",
		X"F8",X"71",X"AE",X"72",X"7D",X"73",X"38",X"74",X"0E",X"16",X"1C",X"32",X"44",X"58",X"70",X"78",
		X"7E",X"8A",X"94",X"A0",X"A6",X"B0",X"63",X"56",X"60",X"6E",X"3C",X"EC",X"4D",X"C0",X"A4",X"0A",
		X"EA",X"6C",X"08",X"00",X"EC",X"F2",X"B0",X"6E",X"3C",X"EC",X"48",X"5A",X"B8",X"66",X"92",X"42",
		X"9A",X"82",X"C3",X"12",X"0E",X"12",X"90",X"4C",X"4D",X"F1",X"A4",X"12",X"2D",X"D2",X"0A",X"64",
		X"C2",X"6C",X"0F",X"66",X"CD",X"82",X"6C",X"9A",X"C3",X"4A",X"85",X"C0",X"A5",X"92",X"BD",X"C2",
		X"B4",X"F0",X"2E",X"12",X"0E",X"26",X"0D",X"D2",X"82",X"4E",X"C0",X"60",X"4E",X"30",X"4D",X"80",
		X"A5",X"92",X"BD",X"C2",X"BB",X"1A",X"4C",X"10",X"0E",X"D8",X"4C",X"82",X"82",X"70",X"C2",X"6C",
		X"0B",X"6E",X"09",X"E6",X"B5",X"92",X"3E",X"00",X"A5",X"92",X"BD",X"C2",X"BE",X"0A",X"B6",X"00",
		X"59",X"62",X"48",X"66",X"D2",X"6D",X"18",X"4E",X"9B",X"64",X"09",X"02",X"3D",X"92",X"43",X"70",
		X"B8",X"00",X"18",X"4E",X"9B",X"64",X"08",X"C2",X"3D",X"92",X"43",X"71",X"20",X"4E",X"9B",X"64",
		X"B8",X"46",X"09",X"EC",X"4A",X"1A",X"C0",X"00",X"3D",X"92",X"43",X"70",X"B8",X"40",X"20",X"56",
		X"2C",X"52",X"0C",X"5A",X"93",X"62",X"CC",X"40",X"34",X"E4",X"CD",X"C2",X"2E",X"03",X"0D",X"17",
		X"1D",X"37",X"4F",X"67",X"7D",X"8B",X"91",X"9D",X"A9",X"B5",X"BB",X"64",X"D2",X"3B",X"2E",X"C2",
		X"6C",X"5A",X"4C",X"93",X"6F",X"BD",X"1A",X"4C",X"12",X"B0",X"40",X"6B",X"2C",X"0A",X"6C",X"5A",
		X"4C",X"93",X"6E",X"0B",X"6E",X"C0",X"52",X"6C",X"92",X"B8",X"50",X"4D",X"82",X"F2",X"58",X"90",
		X"4C",X"4D",X"F0",X"4C",X"80",X"33",X"70",X"C2",X"42",X"5A",X"4C",X"4C",X"82",X"BB",X"52",X"0B",
		X"58",X"B2",X"42",X"6C",X"9A",X"C3",X"4A",X"82",X"64",X"0A",X"5A",X"90",X"00",X"F6",X"6C",X"09",
		X"B2",X"3B",X"2E",X"C1",X"4C",X"4C",X"B6",X"2B",X"20",X"0D",X"A6",X"C1",X"70",X"48",X"50",X"B6",
		X"52",X"3B",X"D2",X"90",X"00",X"DA",X"64",X"90",X"4C",X"C9",X"D8",X"BE",X"0A",X"32",X"42",X"9B",
		X"C2",X"BB",X"1A",X"4C",X"10",X"0A",X"2C",X"CA",X"4E",X"7A",X"65",X"BE",X"0A",X"B6",X"1E",X"94",
		X"D2",X"A2",X"92",X"0A",X"2C",X"CA",X"4E",X"7A",X"65",X"BD",X"1A",X"4C",X"12",X"92",X"13",X"18",
		X"62",X"CA",X"64",X"F2",X"42",X"20",X"6E",X"A3",X"52",X"82",X"40",X"18",X"62",X"CA",X"64",X"F2",
		X"42",X"18",X"6E",X"A3",X"52",X"80",X"00",X"20",X"62",X"CA",X"64",X"F2",X"64",X"08",X"C2",X"BD",
		X"1A",X"4C",X"00",X"7D",X"92",X"43",X"70",X"48",X"40",X"5A",X"60",X"42",X"5A",X"96",X"F2",X"B2",
		X"82",X"56",X"52",X"B0",X"7C",X"DA",X"5A",X"0D",X"E8",X"6A",X"60",X"48",X"00",X"0D",X"17",X"1B",
		X"33",X"43",X"59",X"71",X"7D",X"87",X"93",X"9F",X"AB",X"B1",X"8A",X"5A",X"84",X"12",X"CD",X"82",
		X"B9",X"E6",X"B2",X"40",X"74",X"F2",X"4D",X"83",X"D4",X"F0",X"B2",X"42",X"B9",X"E6",X"B2",X"42",
		X"4D",X"F0",X"0E",X"64",X"0A",X"12",X"B8",X"46",X"10",X"62",X"4B",X"60",X"82",X"72",X"B5",X"C0",
		X"BE",X"A8",X"0A",X"64",X"C5",X"92",X"F0",X"74",X"9D",X"C2",X"6C",X"9A",X"C3",X"4A",X"82",X"6F",
		X"A4",X"F2",X"BD",X"D2",X"F0",X"6C",X"9E",X"0A",X"C2",X"42",X"A4",X"F2",X"B0",X"74",X"9D",X"C2",
		X"6C",X"9A",X"C3",X"4A",X"82",X"6F",X"A4",X"F2",X"BD",X"D2",X"F0",X"6E",X"63",X"52",X"82",X"02",
		X"AE",X"4A",X"92",X"02",X"82",X"70",X"C5",X"92",X"09",X"E6",X"B5",X"92",X"3E",X"13",X"2D",X"28",
		X"CF",X"52",X"B0",X"6E",X"CD",X"82",X"BE",X"0A",X"B6",X"00",X"53",X"64",X"0A",X"12",X"0D",X"0A",
		X"B6",X"1A",X"48",X"00",X"18",X"68",X"6A",X"4E",X"48",X"48",X"0B",X"A6",X"CA",X"72",X"B5",X"C0",
		X"18",X"68",X"6A",X"4E",X"48",X"46",X"0B",X"A6",X"CA",X"72",X"B0",X"00",X"20",X"68",X"6A",X"4E",
		X"4D",X"C2",X"18",X"5C",X"9E",X"52",X"CD",X"80",X"3D",X"92",X"43",X"70",X"B8",X"40",X"20",X"5C",
		X"4E",X"78",X"0C",X"5A",X"93",X"62",X"CC",X"40",X"0D",X"13",X"19",X"33",X"47",X"61",X"6B",X"73",
		X"7D",X"89",X"93",X"9F",X"A5",X"B2",X"4E",X"9D",X"90",X"B8",X"00",X"76",X"56",X"2A",X"26",X"B0",
		X"40",X"BE",X"42",X"A6",X"64",X"C1",X"5C",X"48",X"52",X"BE",X"0A",X"0A",X"64",X"C5",X"92",X"0C",
		X"26",X"B8",X"50",X"6A",X"7C",X"0C",X"52",X"74",X"EC",X"4D",X"C0",X"A4",X"EC",X"0A",X"8A",X"D4",
		X"EC",X"0A",X"64",X"C5",X"92",X"0D",X"F2",X"B8",X"5A",X"93",X"4E",X"69",X"60",X"4D",X"C0",X"9D",
		X"2C",X"6C",X"4A",X"0D",X"A6",X"C1",X"70",X"48",X"68",X"2D",X"8A",X"0D",X"D2",X"82",X"4E",X"3B",
		X"66",X"91",X"6C",X"0C",X"0A",X"0C",X"12",X"C5",X"8B",X"9D",X"2C",X"6C",X"4A",X"0D",X"D8",X"6A",
		X"60",X"40",X"00",X"A6",X"60",X"B9",X"6C",X"0D",X"F0",X"2D",X"B1",X"76",X"52",X"5C",X"C2",X"C2",
		X"6C",X"8B",X"64",X"2A",X"27",X"18",X"54",X"69",X"D8",X"28",X"48",X"0B",X"B2",X"4A",X"E6",X"B8",
		X"00",X"18",X"54",X"69",X"D8",X"28",X"46",X"0B",X"B2",X"4A",X"E7",X"20",X"54",X"69",X"D8",X"2D",
		X"C2",X"18",X"5C",X"CA",X"56",X"98",X"00",X"3D",X"92",X"43",X"70",X"9D",X"C3",X"20",X"5C",X"CA",
		X"56",X"2D",X"C2",X"8B",X"64",X"6C",X"67",X"24",X"73",X"10",X"29",X"8A",X"F0",X"07",X"C0",X"19",
		X"D0",X"22",X"69",X"18",X"A8",X"B9",X"00",X"02",X"C0",X"1A",X"F0",X"1A",X"90",X"2A",X"A9",X"00",
		X"99",X"00",X"02",X"A2",X"E1",X"68",X"68",X"8A",X"6D",X"EF",X"02",X"B0",X"04",X"A9",X"00",X"85",
		X"73",X"8D",X"EF",X"02",X"18",X"60",X"A2",X"80",X"EC",X"EF",X"02",X"90",X"06",X"A2",X"00",X"A0",
		X"1A",X"18",X"60",X"20",X"07",X"75",X"38",X"60",X"A2",X"F8",X"38",X"66",X"71",X"C4",X"72",X"F0",
		X"D4",X"84",X"72",X"0A",X"29",X"86",X"85",X"10",X"30",X"1A",X"F0",X"18",X"B9",X"21",X"02",X"C9",
		X"80",X"6A",X"20",X"62",X"6A",X"99",X"21",X"02",X"B9",X"42",X"02",X"C9",X"80",X"6A",X"20",X"62",
		X"6A",X"99",X"42",X"02",X"A2",X"00",X"20",X"67",X"75",X"A2",X"21",X"98",X"18",X"69",X"21",X"A8",
		X"20",X"67",X"75",X"A2",X"B0",X"D0",X"9E",X"86",X"11",X"B9",X"21",X"02",X"30",X"13",X"BD",X"3A",
		X"02",X"30",X"18",X"20",X"B1",X"75",X"90",X"13",X"A9",X"00",X"38",X"F9",X"21",X"02",X"4C",X"9A",
		X"75",X"BD",X"3A",X"02",X"10",X"05",X"20",X"B1",X"75",X"90",X"ED",X"B9",X"21",X"02",X"24",X"10",
		X"10",X"07",X"C9",X"80",X"6A",X"79",X"21",X"02",X"4A",X"2A",X"20",X"EA",X"68",X"10",X"06",X"C9",
		X"FB",X"90",X"08",X"A9",X"FA",X"C9",X"06",X"B0",X"02",X"A9",X"06",X"A6",X"11",X"9D",X"3A",X"02",
		X"60",X"B9",X"A5",X"02",X"DD",X"BE",X"02",X"B9",X"63",X"02",X"FD",X"7C",X"02",X"60",X"1F",X"C4",
		X"09",X"70",X"2D",X"9A",X"0B",X"64",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"08",X"00",X"00",X"00",X"00",X"16",X"21",X"00",X"00",
		X"00",X"00",X"2F",X"36",X"00",X"00",X"00",X"00",X"3D",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4B",X"52",X"00",X"00",X"00",X"00",X"28",X"21",X"00",X"00",
		X"00",X"00",X"5D",X"64",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"7A",X"85",X"7A",
		X"90",X"A5",X"00",X"00",X"00",X"00",X"90",X"B6",X"D3",X"DE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"C1",X"CC",X"00",X"01",X"04",X"E0",X"03",X"05",X"00",X"00",
		X"01",X"04",X"A8",X"FF",X"05",X"00",X"00",X"01",X"04",X"D0",X"03",X"05",X"00",X"00",X"7F",X"01",
		X"04",X"01",X"10",X"01",X"14",X"FF",X"10",X"00",X"00",X"7F",X"20",X"A2",X"00",X"01",X"00",X"00",
		X"7F",X"01",X"10",X"01",X"20",X"00",X"00",X"01",X"02",X"0C",X"01",X"18",X"00",X"00",X"01",X"10",
		X"A4",X"FF",X"03",X"00",X"00",X"01",X"01",X"04",X"01",X"40",X"00",X"00",X"01",X"10",X"A4",X"FF",
		X"04",X"00",X"00",X"01",X"F0",X"06",X"00",X"02",X"00",X"00",X"0F",X"10",X"A8",X"00",X"01",X"10",
		X"A0",X"00",X"01",X"00",X"00",X"01",X"02",X"50",X"01",X"70",X"00",X"00",X"07",X"10",X"A8",X"00",
		X"01",X"10",X"A0",X"00",X"01",X"00",X"00",X"0C",X"02",X"0A",X"01",X"03",X"04",X"0C",X"FF",X"02",
		X"00",X"00",X"01",X"18",X"A0",X"01",X"05",X"18",X"A5",X"FF",X"05",X"00",X"00",X"18",X"02",X"0A",
		X"01",X"02",X"02",X"0B",X"00",X"02",X"00",X"00",X"10",X"0C",X"21",X"00",X"01",X"0C",X"18",X"00",
		X"01",X"00",X"01",X"02",X"20",X"10",X"FF",X"04",X"30",X"02",X"30",X"00",X"00",X"01",X"30",X"21",
		X"01",X"08",X"00",X"01",X"80",X"84",X"01",X"04",X"30",X"85",X"FF",X"04",X"00",X"00",X"04",X"18",
		X"A5",X"FF",X"04",X"18",X"A1",X"01",X"04",X"00",X"00",X"10",X"0C",X"49",X"00",X"01",X"0C",X"30",
		X"00",X"01",X"00",X"00",X"02",X"C0",X"A4",X"00",X"01",X"00",X"00",X"01",X"01",X"F0",X"01",X"0F",
		X"01",X"FF",X"FF",X"0F",X"00",X"00",X"01",X"1F",X"A2",X"00",X"01",X"00",X"00",X"2C",X"41",X"77",
		X"18",X"90",X"09",X"38",X"B0",X"01",X"18",X"A5",X"22",X"F0",X"F2",X"B8",X"8A",X"48",X"A2",X"07",
		X"90",X"04",X"B5",X"9B",X"D0",X"15",X"B9",X"C8",X"75",X"F0",X"10",X"50",X"02",X"A9",X"00",X"48",
		X"A9",X"00",X"95",X"9B",X"A9",X"80",X"95",X"BB",X"68",X"95",X"9B",X"88",X"CA",X"10",X"E1",X"68",
		X"AA",X"60",X"A2",X"07",X"B4",X"9B",X"F0",X"3A",X"B5",X"BB",X"30",X"41",X"D6",X"AB",X"D0",X"34",
		X"D6",X"B3",X"F0",X"09",X"B5",X"A3",X"18",X"79",X"2A",X"76",X"4C",X"6B",X"77",X"C8",X"C8",X"C8",
		X"C8",X"94",X"9B",X"B9",X"2B",X"76",X"95",X"B3",X"B9",X"29",X"76",X"95",X"A3",X"B9",X"28",X"76",
		X"95",X"AB",X"D0",X"10",X"B4",X"C3",X"D6",X"BB",X"D0",X"E7",X"B4",X"9B",X"C8",X"D0",X"0E",X"A8",
		X"94",X"9B",X"94",X"A3",X"B5",X"A3",X"9D",X"00",X"2C",X"CA",X"10",X"B8",X"60",X"B9",X"28",X"76",
		X"F0",X"ED",X"95",X"BB",X"C8",X"94",X"C3",X"D0",X"C8",X"01",X"E0",X"C0",X"E1",X"E5",X"C3",X"CA",
		X"C3",X"AF",X"C3",X"94",X"C3",X"7F",X"02",X"04",X"04",X"05",X"03",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
