-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu3 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu3 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "3544510691CE55064194935444442188EF09F9D11441A4460739541106526D4C";
    attribute INIT_01 of inst : label is "CAB84635B68686644467DDDD9F568D9C1628E30205D0004A527444538F6460F5";
    attribute INIT_02 of inst : label is "72200565C5488FA58705220656DCD488F95191D95E8F60399997E2D12E242E57";
    attribute INIT_03 of inst : label is "59615223A57152239A214188829181488267B635223A752B888EE64744651A52";
    attribute INIT_04 of inst : label is "6404C41515D204C50D2BADD5A5D515A555A5659440620946949888299C908822";
    attribute INIT_05 of inst : label is "6C5192311B269EA8E284496696A9568FC3A64A8737CB8AD7688BB8515B63690D";
    attribute INIT_06 of inst : label is "22000F8FB2B4216112596D956665E944496CA45A5E5F41115296585D564D045A";
    attribute INIT_07 of inst : label is "8C9999996C07C1B0555557EACACEC96A059E87A9EA7ADC18D452C94E11A734EF";
    attribute INIT_08 of inst : label is "3D866610E24918E94625955466D938F9371F2945614659394D981371E38C548C";
    attribute INIT_09 of inst : label is "1A918895D996620576CC6A674F33AECB10703151E192836DBD068B07ED59F8BD";
    attribute INIT_0A of inst : label is "5DB01A918A95D996628576CC6A674F36F35E979DB4E2E91AE22576E5588D5DB0";
    attribute INIT_0B of inst : label is "A515556926664ADDDD7612501BE88164E2F3697B579DB4E6E91A22A576E558AD";
    attribute INIT_0C of inst : label is "F9BD9526659155551565114584E736E12AA4418155549D101815557425FB1F89";
    attribute INIT_0D of inst : label is "44FA51EEA51E92CA6238FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "0B73DEB41516108DA091528A51E9997F6D92FA84251E6B59A5C6C761916BA323";
    attribute INIT_0F of inst : label is "7FE0452555393939393939393A50FA50FA50FA50F5B15FFFFFFFA533B9384412";
    attribute INIT_10 of inst : label is "ED55555555555530749D24562555571555735C96517B35C94526A1FDFD85287F";
    attribute INIT_11 of inst : label is "623414981546707B5546707B554507B554507B565955555558C9D2772749D241";
    attribute INIT_12 of inst : label is "5C4F6C2786D96A8A89E3AE9992FA4A9A34578D16AFFE6FFE59FEBFBFE3FA4E23";
    attribute INIT_13 of inst : label is "9EB9158EE918F3C912C83A316E399874484693510E78585178D858C5B8E766AA";
    attribute INIT_14 of inst : label is "6994407061535EE6E615DAAA1099D8470CEB6B99D0840ECC1080784745145699";
    attribute INIT_15 of inst : label is "95121AFDE31510E6B6011A6516642E21AA46A11A67861BA11A656886A9286804";
    attribute INIT_16 of inst : label is "0979F41B298ACA580202B44169B67989E2A3E301A68045404689F42910502954";
    attribute INIT_17 of inst : label is "945D9852989924310B89C069492D341A5204679E7463CF3F9D062F6023B8D198";
    attribute INIT_18 of inst : label is "40123611982082042CF3171E1CB33758ACAE2489590626454E11B89A69A16058";
    attribute INIT_19 of inst : label is "2462106BF81C1BB5A289BB56A89B9427C51437154372DD860010991951D00586";
    attribute INIT_1A of inst : label is "4109AF81CBB7E5AA8BB6E56A899B942A8B95A42A489412E50099431A504B9624";
    attribute INIT_1B of inst : label is "02C06C6C6C6C6C6C6318C6318C06451CC3844F3CF62DA0E6A0E6ADB7A870558B";
    attribute INIT_1C of inst : label is "C0602108701C042108701C05B1831B1B1800180C60C4B12C6C1B1B1B1B1B1831";
    attribute INIT_1D of inst : label is "042C018031B000C018312C4B1B1B1B1B12C42C6C018C4B1B1B1B1B1B18C60C42";
    attribute INIT_1E of inst : label is "0310002C6C018318300006C000040000B0000060000300000100008C00000603";
    attribute INIT_1F of inst : label is "FFFFFFFFFDA170BDAF721C8721C8721C8721C8721C8721C8721C8721C8721C84";
    attribute INIT_20 of inst : label is "61CD18F2003761C1580C2F1D0C608A40186593CF3440C2FFFFFFFFFBAB87AC4B";
    attribute INIT_21 of inst : label is "6862A6D36DA3C54135E5112F94541424E49CE3E242B4CE4A09112E1BD9870E07";
    attribute INIT_22 of inst : label is "0212DA4C44BE760210D145B04E6D051CEC6DCCDA90E2FE2581981982988C6A61";
    attribute INIT_23 of inst : label is "080159666BCF2A60B00002022002122751127511C447111F446AC449C4B513C6";
    attribute INIT_24 of inst : label is "490F36693CAA1B96890F36A9006A19299243CD9A422A8644105771F83002DC95";
    attribute INIT_25 of inst : label is "6429B5E1C50B94EE446D0E10B6808B253BCC9A3F9044E96A243CDAA4D1A864AA";
    attribute INIT_26 of inst : label is "8B1BBA303FEE2279E3CEE28CFB9889168B04A925DB092716063C687046F5425E";
    attribute INIT_27 of inst : label is "B989EA2179B5AA8789102330009FFD000AAAAAAD9D033AA8100580C2F3C2A137";
    attribute INIT_28 of inst : label is "65547DE47FFE26C0E4298E2C2728A7222D541A5360435420E10B0550FEFFCF07";
    attribute INIT_29 of inst : label is "5A738B06AE060D87242E0D841041BABC741C31B6D86CC6EC66C4B011EFF5545D";
    attribute INIT_2A of inst : label is "0B0644D7491406B47080B0E41A514A918AD1CDBBBEDD67B499A6598ED9B8FAEB";
    attribute INIT_2B of inst : label is "00730330C40796262B06BE04031000754E519511519B98D9D052450106847080";
    attribute INIT_2C of inst : label is "16A499455DC626163362A6C1BCAA62F4A053507A054D5595D2C0CC301C31012C";
    attribute INIT_2D of inst : label is "601B63169898AC1AF814EB36AF755D4D555D575355096AAA24446ADD11B65165";
    attribute INIT_2E of inst : label is "3DC7F61FD45F417FA38B100BEAE9ECC0CCCCC705F60B609774B3033331C070DF";
    attribute INIT_2F of inst : label is "00000002A940FFA9403FA55D1E615DE62B06E812C58B1D08F36C2DAC1A36FA6D";
    attribute INIT_30 of inst : label is "BEDACC648B6F3CF3CF3C8BC191918700A1A8084A1546400080050DA68CEBBE80";
    attribute INIT_31 of inst : label is "2C54D8536207361CD88C54D8536207361CD8AC1804B86D999951FA6C46F68437";
    attribute INIT_32 of inst : label is "1F3338BCCE3FAECEA8B612D04B62832F6018104F6EAEA7BED8063893A838B390";
    attribute INIT_33 of inst : label is "6102612CFA6D29B6842360A6529A60D46626FFA652CFA6261FA6D29A0C546CCE";
    attribute INIT_34 of inst : label is "652CFA6D20FA6529A60D46623FA6D20FA652DFA612CFA6129A60D4618DB3E540";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF61B4264DA61A1101B402CFA";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "109423FD6161E996911670013EE7A6447BD3D8280B04E1AFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "C840C8504444478378EC55C8F91062F800000000000000000000000013BCA1C5";
    attribute INIT_39 of inst : label is "3FA5DCE0F297F383BA5DCE0E2977F834A5CFE0D297FF834A5EFE0DE977F83440";
    attribute INIT_3A of inst : label is "B725EB8695F620E92136B0667C06004E9021154D7F791252D43A5DCE0C297B38";
    attribute INIT_3B of inst : label is "8E69502F955DB00431A2E0F5DB00E68C5E50D13C104509818374A668E5590290";
    attribute INIT_3C of inst : label is "158509000000195C8824596EC52A74034EA4ADD946550E4A05CE8C170A390541";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC8D44168F28966917CF0DC7CE5";
    attribute INIT_3E of inst : label is "5E818851B2644A1A13063CF3391A558923411709341041A853FFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFF286BD991581C55859D47185314E64048674001118585185985314E";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "67888A2BEF998619C4236C58888B0000C24A0D62228AFB090E66186F10899132";
    attribute INIT_01 of inst : label is "1D7572814485B4DAC8F9AAAA024893A015089437DFFC491F6288FC5250A811BC";
    attribute INIT_02 of inst : label is "F4E6E4675B5395E1AF7F4E63C6B5F53961BAB6B243074C622221B9360B983445";
    attribute INIT_03 of inst : label is "49D6C4E575C6E4E50E6B1F9398DB5F53983DAD7C4E526D42939486EADBC998F5";
    attribute INIT_04 of inst : label is "C472B04A398BB2B848B2B7AEAC0A38D90939390BD7EC4266317939993575398C";
    attribute INIT_05 of inst : label is "D387450656F362852CD8C0D0C3C4D24106566189DD13A27A998399FB72D7E39F";
    attribute INIT_06 of inst : label is "4E6AA2A297AD4FC63034FF3B88838898C0D3810C083B0631BC0D0D090D7018CD";
    attribute INIT_07 of inst : label is "062222097383A0EBAAAA8E9730393004536398EE3A8EEFF1B945BC8D605E7520";
    attribute INIT_08 of inst : label is "39F6AB05D77E1F2096C2530A79BA252548AF50A08081A63683AFA34E92505606";
    attribute INIT_09 of inst : label is "1536E2A7F07DB899FC0C54CA7B7BC8A8DD4DDD6390A16B4D35549A11884415A6";
    attribute INIT_0A of inst : label is "7F001536E2A7F07DB899FC0C54CA6B67B647C74378D6B20578B9FC5F6E2E7F00";
    attribute INIT_0B of inst : label is "196AAA8948888EAAAA7E13A232104148D637491E874378D4B205F8B9FC5F6E2E";
    attribute INIT_0C of inst : label is "F7BDAE2B92ECB9E609926F9AD2AF1494B12482FAAAA8262230AAAABD09271807";
    attribute INIT_0D of inst : label is "5290A1B54A1BCB674F75FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "20F4F8D74A39B110D361452CA1B22219D3209D4C4A1B34C01791BC0E2F92A4E0";
    attribute INIT_0F of inst : label is "91F00CD75595403FEA95403FE800FFFFAAAA5555000555555555554400407820";
    attribute INIT_10 of inst : label is "131DD57754000008FE3F3805315555F800D0E4FB33050E4FA331526644DCD499";
    attribute INIT_11 of inst : label is "E12C0E3C081CD012581CD012581E012581E012587600CC03342F7BDCBDEF7380";
    attribute INIT_12 of inst : label is "898E9840470807CD3833D622219E0F7E308E8C220FFE0FFE4BFEFFAFEFFAA292";
    attribute INIT_13 of inst : label is "3CEA0CD0987977522339654149263C488D8140279094ACAF3A3CAD05249860FF";
    attribute INIT_14 of inst : label is "8826D6C6C7C7CC62A37E3F35B1E35B9C09D3CE352CF8A190106EF058B82F8335";
    attribute INIT_15 of inst : label is "82E290AFCEB6F90A83C4A20984C54C4A309094A30BA33194A309A528828CC712";
    attribute INIT_16 of inst : label is "D4F3A80C0715454E2F895400B3E8E3F38FCE9411455057804D33B81500244278";
    attribute INIT_17 of inst : label is "22A022AC236635060651045D04FC1015E004D33B8BE5DD6C6A00D0D75DADE075";
    attribute INIT_18 of inst : label is "E4DF6EC6B1F7DC71F6B980F4AFDAC071545B7B138A38D99D8D606DBCDED412A4";
    attribute INIT_19 of inst : label is "D4E3E202941512C51EDD2E51A5D2D5D69AF90D4790D7931C71C6A205E431371A";
    attribute INIT_1A of inst : label is "82820A4152C7981ED2E7581E5E62D4DE52D798DE1E6C679B15F6C579B112D798";
    attribute INIT_1B of inst : label is "03C00156ABFC0156A2FCC00546068E338214B775AE3911756171EC4FD8D35F8D";
    attribute INIT_1C of inst : label is "B0F010060DC070180405C272AFC30055A80000015068AF3C0055AAFF0055A82F";
    attribute INIT_1D of inst : label is "14140A802FF000B03C300145AAFF0055A2BC3C0005468AFF0055AAFF00150682";
    attribute INIT_1E of inst : label is "03000001540A82FC3000000000140000580000A0000200000F0000CC00000000";
    attribute INIT_1F of inst : label is "FFFFFFFFFDB6CB186F864090E429064090E429064090E429064090E429064090";
    attribute INIT_20 of inst : label is "E18928E14524E18971241758717452716BCD6DDD678821FFFFFFFFF08E8638C2";
    attribute INIT_21 of inst : label is "000846A32010651A02027708080B0A1B36E7107EF56841460D73081ED3864E24";
    attribute INIT_22 of inst : label is "FF55855552426EC3600000604567DF7D04D3D04D41D3544B5575675771A45408";
    attribute INIT_23 of inst : label is "0400233BB1DD51BDD5D649649649549095490D5415509541552415351501541E";
    attribute INIT_24 of inst : label is "20334D20150003802033412039000020080CD3480D40003DFBDFE088200228EE";
    attribute INIT_25 of inst : label is "A810B0126184E0A0981F12605E054DF408D1489503904D3080CD04806400008C";
    attribute INIT_26 of inst : label is "45844D0415DEB48510651241537AD23445B5DA3CD8A42F4DA613049A69820C20";
    attribute INIT_27 of inst : label is "6C95D3254C95BE777EC5E7C7F42AA9AAA5555559921D7480D00712417751FBB4";
    attribute INIT_28 of inst : label is "D34DE34AFFFD0FAFC20FCF8435B6C4BCB540C70214414BD070264540A2FFCA77";
    attribute INIT_29 of inst : label is "4ACCE4595814745CF458344000002564F8A6455003FC6A815FC0AC839FF38E34";
    attribute INIT_2A of inst : label is "044940C73CF3B4A5C400449712171A171217133D3873FD668D237228323614D5";
    attribute INIT_2B of inst : label is "00403C03C444BF5D44496436E3188445334454454411514543810401A495C400";
    attribute INIT_2C of inst : label is "FAA8A4B2473EDF7D714101125A556616B1C7D05BF71FFF130F3F000010F111A0";
    attribute INIT_2D of inst : label is "C013C01A3D75112590D336515945131FFF5144C7DF113154346B8E9DAE5EE092";
    attribute INIT_2E of inst : label is "03140C503140C540875CCF4194F9200F0003C59B3CF3C116C3C03C0031005973";
    attribute INIT_2F of inst : label is "00000002AAAA55555540000D719CFF3BC45990DB312CC71345184F1164116541";
    attribute INIT_30 of inst : label is "38F119974917757757756F5F2F206C966320A8C8189C8009800F133D1093D940";
    attribute INIT_31 of inst : label is "33253D94D4FB4F6D350C693DA4D4084F61351126CCAA2F2222FE65732E0EF84C";
    attribute INIT_32 of inst : label is "351114D445355CC6698F6239A8D4718E7EFC715F4D351C38F044658669648650";
    attribute INIT_33 of inst : label is "CB1310DC671CDC60B1E7C071C1C7146171E1F6718DC671D1067141C546217445";
    attribute INIT_34 of inst : label is "14DC6714D067181C5146171D36710D06710DC6710DC6714DC4146170707194C4";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF70401A9F314287132C4DC67";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "03533725D4D795D75C450FF30975D43115F0B5D40137D1FFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "3333FFFF7777752FEF4827D1CF23535400000000000000000000000010B5104D";
    attribute INIT_39 of inst : label is "F326CF4BCC9B3D2F326CF4BCC9B7D2F326DF4BCC9B3D2F326CF4BCC9B3D2F377";
    attribute INIT_3A of inst : label is "BD3B94E5352ED07630316457900784694323268620FD41C090B26CF4BDC9B3D2";
    attribute INIT_3B of inst : label is "7041C4D81556C806015D5061EC8835443A7DA010000537116968CF98972C0148";
    attribute INIT_3C of inst : label is "82023600000044525C7D45539C51B6EF6374F91C47DC704D57D1701F45C1F711";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8D4000418457B009DD522BDC2";
    attribute INIT_3E of inst : label is "833037C56F79852F2FDE5DD68A058E355713504C20830CE8C3FFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFF683FDEE209A28B5A70A5BCA41499B79A43DDDDA2CA4AB5AFCA4149";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "CD044D36D7A24125CC99D3E0444520886F8D3B41134DB56B0E890497326B4F15";
    attribute INIT_01 of inst : label is "F2DAF2CBF84849F485A51111E0F0E3D4060EB30A672F8EB6C0445C1ACC46B24A";
    attribute INIT_02 of inst : label is "FEC88837F7FB24A0EFEFEC8243FFFFB262E1A16DE18489E1111B0B2140780782";
    attribute INIT_03 of inst : label is "A6CECEC92BCFCEC9CA13333B20A7373B23266CECEC91BCC93B278A8486B7B0FC";
    attribute INIT_04 of inst : label is "7C6813890621A81D8210EF592CC906F717171714CCC8C9EC3333B2067373B238";
    attribute INIT_05 of inst : label is "66D86330287BD3CA34E80AF861BEDBC338ACE2F48F21C2947691FE422E8CAE32";
    attribute INIT_06 of inst : label is "ECBFF3F3D28CD8CE02BED2E6447B18280AF0C28783B13A0233AF84836F24E82F";
    attribute INIT_07 of inst : label is "811111ADF5CB32CD55556C2B51C2598CABD0D4390D43D23330AF1D67D8EEBA3E";
    attribute INIT_08 of inst : label is "93DD47E832943D2258892625B67DACCB24D78353436B719F0BDDC1BD2ACC1D81";
    attribute INIT_09 of inst : label is "5A79D7522A8C75D48A4F69E637FCEA9546D4E3A023DAD7AD8C20C1392A4E6C55";
    attribute INIT_0A of inst : label is "22905A79D5522A8C75548A4F69E637F37FE5A6E4F670794EF5E48AA31D7D2290";
    attribute INIT_0B of inst : label is "B715554204447A1111EBE3C3E8E8C5D670FF0F9766E4F670794EF5648AA31D5D";
    attribute INIT_0C of inst : label is "F3FF992759D267151555D077F81FFABE193D01DD55549813E0D5554824CBD3AC";
    attribute INIT_0D of inst : label is "8B1E8292E829610D89DAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "38CD2E118906738E3AD063BE829111B032D40BA8E8298C9A7EFB3B3C1700D4B3";
    attribute INIT_0F of inst : label is "7BF256091BAAAA9555555540015500000000000000000000000000000000D012";
    attribute INIT_10 of inst : label is "056E64B9924E4F6028CA3C20571B188392765CD1959365CD095935EDECD60D7B";
    attribute INIT_11 of inst : label is "7B05240E22D5A27AE2D5A27AE2D507AE2D527AE24C1A6C69B984A02A0280A3C2";
    attribute INIT_12 of inst : label is "046404EAE92DAD671E997F111A3BA69F3C76CF1E9FFE9FFE58FE3F8FE3F89BB0";
    attribute INIT_13 of inst : label is "A60C1A8EB0A6492C13528A306BAD84904D638CD332505057972058C1AEB4BA65";
    attribute INIT_14 of inst : label is "449DCFCECCCCB6D1D2213D8E2392864B403CA08FC4F0CE0C94F198D4430F7A8F";
    attribute INIT_15 of inst : label is "89C52EC36C6173254DBCD127C888E7CD224C8CD22573EA8CD2272B3449CFA2F3";
    attribute INIT_16 of inst : label is "1D9B3037AD65DBCF33CE9CC378760B5B2D6C19018AE26B005FDB363B30D3C9E5";
    attribute INIT_17 of inst : label is "9350935899D9013D8C62406ECB3F2C9AC305FDB3719924839C0E737833C6D8DE";
    attribute INIT_18 of inst : label is "1A538C184A18E086553505555D5405D65DB1B7E04D3676586758C626FD497354";
    attribute INIT_19 of inst : label is "BF93C33A18912A493112A49F552A49BDE84AB088AB0A0C60861B794F28CA94E1";
    attribute INIT_1A of inst : label is "01C9E8891A4875311A48B5F553DA49B95A4835BD13D38434E13D38434E1A48F5";
    attribute INIT_1B of inst : label is "0283FFFFFFFC0000000015154509EBA2103F14920893F1CB11C710D8B0B97A4F";
    attribute INIT_1C of inst : label is "F0F069180B52C065190353C15541AAAAA80000000000000154555555AAAAA82A";
    attribute INIT_1D of inst : label is "68295A802AA000A0282F3FCFFFFF00000000015455554555AAAAAAAAFCFF0FC3";
    attribute INIT_1E of inst : label is "0300000000001400055555555555555555515555455555155555554555552A56";
    attribute INIT_1F of inst : label is "FFFFFFFFFBEFBEFBEF9785A1184D124451F0781D07E1A8661B4691545C160540";
    attribute INIT_20 of inst : label is "CA297E47DAA4CA29D69D34B786B9E126B4CBC5248F0DEFFFFFFFFFF5D1284690";
    attribute INIT_21 of inst : label is "E0E9ECC3CDF0E1410D0D2240363536357E8D50F26A80EFD3863A43A4E3281FA4";
    attribute INIT_22 of inst : label is "435A170D65CCA943C0F3CF825B0DE69E0D75E0D791B05F25E6DE5DE4D65D3CE4";
    attribute INIT_23 of inst : label is "8C08D6177924AA5649E69B69F69F5933A5933A58E963A58E964CD64CD63258F9";
    attribute INIT_24 of inst : label is "09959F39AF2A3B4609959F399B2839B1826567CE65CA0EACBACC840500136459";
    attribute INIT_25 of inst : label is "563E7DF0E59C5642563635D8C885C199B164CE1FD9368A1826567CE68CA4E6C6";
    attribute INIT_26 of inst : label is "C39FDF303F322251F0E3F8CC7CC88987C3853C0AE38DB79784397C3863056492";
    attribute INIT_27 of inst : label is "C9513A546A59E554D89DBDAE8C97748881393933FC08CC88F00D69D3492A657B";
    attribute INIT_28 of inst : label is "451410457FFC1451D4151D605D16491596CCB732E04BF150F3380730A1000A74";
    attribute INIT_29 of inst : label is "6EA5C69FA206B5FA74A235CC30C38E84B80A800A815655555014005A5FF51451";
    attribute INIT_2A of inst : label is "069FCCE7CF3CF878BC8069FD212231223522329593F2DDC7CD733DB23DAF1E79";
    attribute INIT_2B of inst : label is "02620223E4075FCFE69F863F339CC04B174A84A84A8DD65FF0F3CF09F878BC80";
    attribute INIT_2C of inst : label is "06649649C6995FCFFFA3B1A7D00084DF50CCA0750332FFFE8780882098F10158";
    attribute INIT_2D of inst : label is "A01CA019FF3F9A7E18F17597A1CB2232FFB2C88CA3333C03ABB77122DD951155";
    attribute INIT_2E of inst : label is "323CC8F323CC8ECC8DAD4E8D2A1A58808888E52BCA0CA01FA1E202223982527C";
    attribute INIT_2F of inst : label is "00000002C586B16CAC5B6B17AA6CD277669F28FB532D42317970729A7E174ACF";
    attribute INIT_30 of inst : label is "B329A1FB8D7492492492812F9E94CA5B1E18C786164E4004C00232A38EBB5280";
    attribute INIT_31 of inst : label is "35162F58BE048BD22F8C522F48BE048BD22F9A7CBB48121111424AF50A69D48B";
    attribute INIT_32 of inst : label is "1C000470011C6FCD75CBD3234CBE732CF4E4338F6BAB1BB328044844844944B0";
    attribute INIT_33 of inst : label is "927B535ECB5F2D7C7C9D90B5F2D7E0DAF54DDCB535ECB54D2CB532D60CDAF001";
    attribute INIT_34 of inst : label is "5F5ECB5F52CB5F2D7E0DAF551CB5352CB535ECB535ECB532D4E0DAF35F732CAE";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF37C227675F1F2BA49E5CCB";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "39F169C779797659249BFFFE41964B126D241E5C0F953A6FFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "9D1559D11111115351506DE13C21B07800000000000000000000000035D2F3E5";
    attribute INIT_39 of inst : label is "3385CD54C6173553385CD54C6173D53185CF54C6173D53185CF54CE173D53115";
    attribute INIT_3A of inst : label is "4933B3A3776952FC333E806E0427007E93302F03B341065541B85CD54C617355";
    attribute INIT_3B of inst : label is "CC9559F32A78DC2701A512C78DCC36805BDEC30C30C19D64D7D0CA44B31D0B84";
    attribute INIT_3C of inst : label is "0D0D9D0000006C8EA69E6C8D25AA7F30B7C9526591258C9755E6CD5793320564";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6DCC37C39E9F7835248935E0D";
    attribute INIT_3E of inst : label is "61838E8E87F56B86C5A99248358E718F092CB3031C70C77C33FFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFF3E9BFD41041343853249705306B65706BC8CCF810505385305306B";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "9BBFCF3F3C2DC30C4C3672BBFFFDF3FC308F2EEFF3CFCFD900B70C3130D9CA3C";
    attribute INIT_01 of inst : label is "324293C640203070E0E188885DB9A1CD0075127861129E6FE501800448111685";
    attribute INIT_02 of inst : label is "4C09C1913130245644C4C09119131302503430349F1400D000064D3084D53413";
    attribute INIT_03 of inst : label is "005C5C09145C5C096545757024557570251115D5C09155D2702541D1C0D2A04C";
    attribute INIT_04 of inst : label is "0AC774870DDFC770ADF57D4C30870D9E3E2E2E3C4C40C3A8171702451717025C";
    attribute INIT_05 of inst : label is "0008DD2107C6765E41673197DFE986437B18A640042676E10E66462310CC5331";
    attribute INIT_06 of inst : label is "C09555455144C04DCC65B1B300164DA73194567E756749CD19197F76990D2719";
    attribute INIT_07 of inst : label is "3C0000188FF67D9E222219C4F7DCF375267751D4751D80131419F015C4508E6D";
    attribute INIT_08 of inst : label is "56391018E17E6330E003830D0D1C44B62CF1A1D1E1D1F85791C3E5F0D448083C";
    attribute INIT_09 of inst : label is "0110084313460210C4DF04434BCCCDBBDEBDB41CCCC44F1C7DE55E3759D9C9A4";
    attribute INIT_0A of inst : label is "313401103A4313460E90C4DF04436BD6BD9FDC9EA15780854210C49100883134";
    attribute INIT_0B of inst : label is "9EE222200000054444BC84EFD094408157FC567F1C9EA15580854E90C49103A8";
    attribute INIT_0C of inst : label is "F47E84E330C012C4C130C3333747F98DF15BBF3E22203EF7DDE222040CB7C264";
    attribute INIT_0D of inst : label is "4664F0C64F0C5F6400C2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_0E of inst : label is "3C4F15D7870C1309D4701DF0F0C00065D348594CCF0C7471D3364C1E0F8FC022";
    attribute INIT_0F of inst : label is "11C0380FFF00000000000000000000000000000000000000000000000000BB7F";
    attribute INIT_10 of inst : label is "0D3FFFFFFFFFFF07DDB70000F3FFFDFFFFF0C4743E030C4743E0304444380C11";
    attribute INIT_11 of inst : label is "F13E0D750FD5E215FFD5E015FFD4215FFD4015FCF7FFFFFFFC1F77DC7DDF7000";
    attribute INIT_12 of inst : label is "681568C75737769535F5C50004457F0D75135D440FFC0FFC00FC3F0FC3F0C313";
    attribute INIT_13 of inst : label is "F51EFCC9148628EE7CF5B12011474C39F111407170EC383103343C80451CD7FA";
    attribute INIT_14 of inst : label is "C4394C4C4C4C44818130D2453343420CC4E45146ED3BC9C80C70D39001C40346";
    attribute INIT_15 of inst : label is "C3E105115130170F072CF10EC0C0CCCF10C4CCF10F33D3CCF10E7F3C43CF40B3";
    attribute INIT_16 of inst : label is "54D47B124560F98370DD6841C4F114D453515B4000E0239135546116107BC390";
    attribute INIT_17 of inst : label is "33EC33EC3577332C4560D0035D0D7405E5135144FB18A3B67EC55249545A8452";
    attribute INIT_18 of inst : label is "690784681679E79A00300E000C000D960F968C60CF0D5DCC15445AB9130B93E4";
    attribute INIT_19 of inst : label is "9BE4EF15640305C390305C310305C399EEDA2681A26BC9659E6B3086689A4120";
    attribute INIT_1A of inst : label is "BFC3554035C1DF9035C1DF103575C39035C1DF9034758D1D634758DDD635C11F";
    attribute INIT_1B of inst : label is "000000000001555551545515450CC750A13BB28ECC56A0D500D5064D90342F93";
    attribute INIT_1C of inst : label is "A0A0982445415898244941595541555554000000000000000000000000000000";
    attribute INIT_1D of inst : label is "BC3EAFC03FF00050141515455555AAAAA2A82AA8AAAA8AAAAAAAAAAAA8AA0A82";
    attribute INIT_1E of inst : label is "02F0003FFC0FEBFC3AAAEFEAAABEAAAAFEA2AAFA8AABAA2AAFAAAACEAAAA3FAB";
    attribute INIT_1F of inst : label is "FFFFFFFFFAAAAAAAAF8E6398E6398E6398A6298A6298A6298A6298A6298A6298";
    attribute INIT_20 of inst : label is "455445571A504554960F92A69A09E4068046ECA3BBBC91FFFFFFFFF452154861";
    attribute INIT_21 of inst : label is "787478EF49A0D043070731841C1D1D1FCAE7F0C34930D5958D11855EC1159150";
    attribute INIT_22 of inst : label is "C049F10D2E483EFCE51451703D0DA5920FDD20FD1553490D25525525560F9074";
    attribute INIT_23 of inst : label is "4400732CCCA39DDA5924BD4BD4BD4B9204B920488122048812C492C4922048BE";
    attribute INIT_24 of inst : label is "0DC6993DF30C1C0F0DC6993DCB0D1DD3C371A64F73C3870104346842101148B4";
    attribute INIT_25 of inst : label is "D1143520D044B780D113B4C44C164DD5F1A74F4A5C37C52C371A64F7CC30774B";
    attribute INIT_26 of inst : label is "8344B9202AE310FC20D12648278C436283419ECCC245D4B5403B683411CF7030";
    attribute INIT_27 of inst : label is "8438E10E043410C3941C0C0C0C3940A503EA9542EEC0F8E3200960F928E4F230";
    attribute INIT_28 of inst : label is "000000003FFC3C00C0340C00FB3FC337F4851C145003B9F2C1770214B0554BE3";
    attribute INIT_29 of inst : label is "67CF04BD4CC4877CC49CC7471C71453A3000000000000000000202000FF00000";
    attribute INIT_2A of inst : label is "04B995F04104C000CC004BDB000330033003314C45D101B54150143814471916";
    attribute INIT_2B of inst : label is "502642ECF10004C4C4BD78CB37CFD0023C79979979959E76141C5140C000CC00";
    attribute INIT_2C of inst : label is "33238C008F3EC4C4FF91112F6F004CAB144C51310131006B0C80BB64093C4009";
    attribute INIT_2D of inst : label is "444444C0131312F5E323C79D4E820331006080CC513E04021F0111B0046CCC30";
    attribute INIT_2E of inst : label is "23388CE23388CD88CC23C08EC538C990BBB8F16D0404440AC32642EE7C901610";
    attribute INIT_2F of inst : label is "000000025264949225244942F1C471CCC4BDD328F223C33F69DCD112F4DDB18A";
    attribute INIT_30 of inst : label is "45112FD47DD28E28E28E0CED0F087C6B1D13C744D00400057FF3316A0914EC40";
    attribute INIT_31 of inst : label is "CF123348CC048CD2331F123348CCF48CD23312F5F76511000001B18F3CFE358C";
    attribute INIT_32 of inst : label is "0CCCCC33330CDFFD544CDD3764CCF3518CF5134F1162CC451100F40F40F40F6F";
    attribute INIT_33 of inst : label is "63FCB5FFF4B112C4040C6F4B1D2C50D68BD7FF4B5FFF4BD70F4B5D2D0D568333";
    attribute INIT_34 of inst : label is "B1FFF4B1F0F4B1D2C50D68BF0F4B5F0F4B5FFF4B5FFF4B512D50D681F1FFD8FF";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81C7D3318B1013BD8FFFFF4";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "146348BA49491CF305B10AAD873CC116C6185254034115FFFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "99DDDDD1999998030000D92320D55364000000000000000000000000254EA0D0";
    attribute INIT_39 of inst : label is "3300CC00C0033003300CC00C0033C03000CF00C0033C03000CF00CC033C03199";
    attribute INIT_3A of inst : label is "46B1E2D1E2FEF0CEC175700BBD0010351CFCDBBF12000F0003F00CC00C003300";
    attribute INIT_3B of inst : label is "48147B920F2E3D034C1F30FAE3FD30739D9AE1491440456E43BACE03E1814140";
    attribute INIT_3C of inst : label is "078747000000F4082386E408A39DFB313D53B4DD3B47883951AD4946B92051EE";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF108716834508CE1CA38B3C607";
    attribute INIT_3E of inst : label is "DF0144CD7C8D115FED618A3B6445C0464960A2114514513517FFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFFFF553FE3E70033C14310D21432011DCF85106AAAE783831431432011";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
