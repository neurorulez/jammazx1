-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GAL_FIR is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GAL_FIR is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "588552E96981EFA5D6A0EC4DDE65766C0563812E830944010D0D1100066709A6";
    attribute INIT_01 of inst : label is "56298A03D5EFE3EED97416D80902F8B33C5D02FEC4BFB42E46D5A9C57FD2BA05";
    attribute INIT_02 of inst : label is "11F8207EF9CA1AFF9F8128EBF28FBCD3A0BF16E9AAFC9374F028805EAF3EB667";
    attribute INIT_03 of inst : label is "D41ABAAED4BBA8CC52F5F24FBCAE6CA58AE384E274A0A16C836142AECEFBEA73";
    attribute INIT_04 of inst : label is "356F94FB9924F3609EE9990367972EE54D10D8669E729AEFC8C2471B6BD881E5";
    attribute INIT_05 of inst : label is "32E4F4B1E6E66BBB9E0D297616AD9E2BD23AA43B43578A3A852EB0550A11A0D6";
    attribute INIT_06 of inst : label is "0BE72F93A40705A8AC6800DB6A4D2DF323B722CA4A3A694CC0CC886BB07B7DF9";
    attribute INIT_07 of inst : label is "11C6535CCE0A74517260EB76621142DE73141FE0EE738794FCD3E9888B39B7DD";
    attribute INIT_08 of inst : label is "6DDA99282AA319CB4657D7A04980E2A2EAC6A0778AFD9923A82CAD25A1986AF8";
    attribute INIT_09 of inst : label is "DCFA72CBD0ED6854C56DBB7C04988809EE0B7D80B9196912CEC9E6F6FC720257";
    attribute INIT_0A of inst : label is "9040C874DDB2000F9794689CC1115D6F24629904F6EC8CCC557918FABAED3E44";
    attribute INIT_0B of inst : label is "90592B8FF6648992227BDEB5490C3306E7A138AD804AA21C566BD19AA53090AF";
    attribute INIT_0C of inst : label is "94533F03DCBFD18B4E8F1592BA80D3E4CE29A7881607D43ECFBD45747B407CBE";
    attribute INIT_0D of inst : label is "7ED4B7A65EB96284E2B1FB3A3C792A261E3754B0715878D45E9F810FE39C2B71";
    attribute INIT_0E of inst : label is "9D5C35EE6AA7E861D4E490BAB0350DE8D16EF8810F82FA330F949B1C74720AB3";
    attribute INIT_0F of inst : label is "ACDB0735AEA73F1EE614765A516A0258332A15405F5AE1F9FF1621A95742729D";
    attribute INIT_10 of inst : label is "67F927AFDD2648D0302996D692F47CCCCC152F5D3FAD8BF9263584A1D531D369";
    attribute INIT_11 of inst : label is "A6515B7628C79FA94E4AD19A581EE8174C63332B8F722BA5780B3D84C6FF42EB";
    attribute INIT_12 of inst : label is "6C7C22E6D8F7CF911B636EA3C3A282E1E6A3CBFD6241A126556B47EF8E1EDDF9";
    attribute INIT_13 of inst : label is "2F3CC6332B2B2FECFECEFBDBFED6D61C4EB06D7EC1A62A2446FDB1171B2871A8";
    attribute INIT_14 of inst : label is "5E62355DB95BA35CC2BC5E723C35BEED91D423AB6DA348FC63B4D6DBEC6C6B86";
    attribute INIT_15 of inst : label is "7F9CD99AC3A998DD21A21F2E0A22BAC02D3F0EEC305714EE0DE4DA4CD616B83A";
    attribute INIT_16 of inst : label is "1E7F1C1819268726758508F0376EC928A1DDFE3FECB82BF78E2602899D4056CB";
    attribute INIT_17 of inst : label is "4433A34FB4043B7D838D31D7987D9FE3EB4723141E8ACB58963DC14D5B9FE0E0";
    attribute INIT_18 of inst : label is "297C24664DA52671DABF84F1F4654444091A0240BF500836F6AE51A5400125E2";
    attribute INIT_19 of inst : label is "E24A9D49CCAD3DB052DE013540A133921AC16860866DA736588AAD3497CD5CF3";
    attribute INIT_1A of inst : label is "005556DC20D7FFE5212F694C0AACDBFABAE779560200B67B73FD4DA1A36B7895";
    attribute INIT_1B of inst : label is "56EFC33E485819D2E9CEB61877086187ACE92A760F730F446243F7B48F5D2C1C";
    attribute INIT_1C of inst : label is "E5E077C380BFE2D8F9F11F9448E022669B4026A863171004686D474DEECCA291";
    attribute INIT_1D of inst : label is "7F40C3F06EEF6565BCAC924320A1C367A8EF96E02D1740016945E3ECF9584662";
    attribute INIT_1E of inst : label is "718150F3E88DA66744D6665B9DEB54F420576B6800C486917B3DCE351D9F5AE0";
    attribute INIT_1F of inst : label is "888B7522671BFA3EA965018CE6900875B0203905C8CA713FC7B6ABE97F092875";
    attribute INIT_20 of inst : label is "B69852F6E9BDD19B0038EBBDBEEB7B36FAE6C74119E7453CE302F17805A51EAD";
    attribute INIT_21 of inst : label is "3AFED5E24D1FAB979BFDEA51AC482A6BBFB33A92C12A26492DE55411FABD6D71";
    attribute INIT_22 of inst : label is "DC5410D51E3F4C138B7FEA0ED02C42684C288311C0D4A2737BF0E1024E2E6E52";
    attribute INIT_23 of inst : label is "30993FB7F50CC3B841C6C571E74F77A90B4C8354B0F991FB7FFA0B48C580AFF2";
    attribute INIT_24 of inst : label is "7A3EF2B6104C447696914C02CA6DE401FC872E2BC5A03B220120D709B5EC6B37";
    attribute INIT_25 of inst : label is "DC60E13434E3363043573CB2974528F4EC396970694679BD46C70E8EFB26C4BF";
    attribute INIT_26 of inst : label is "B35F9E9126B0F0A78CE7B8DC84BF435283F9D8A481C627235F440F7FB33D0281";
    attribute INIT_27 of inst : label is "53B79F4E0D283725D928E32D422167AE52D606C975E95D9DD9CF5402BDF3E433";
    attribute INIT_28 of inst : label is "B624E88F5E1C24F6E4B2CAF95467DC337211B26D3CA48C26178F1EDF27839E56";
    attribute INIT_29 of inst : label is "9E647AFCA9179241457518F8C18768650D893A7D17D824F5C29EC0392CCEFAB7";
    attribute INIT_2A of inst : label is "79C134E5F03C60E300AA9A4A994C3A044CCCF9E8FE885429145198F53060C7A0";
    attribute INIT_2B of inst : label is "135343398A9F235084CECF20D762F860D832571C4F7F48284579BAAA260D7793";
    attribute INIT_2C of inst : label is "B093429F65E5ECFC35B8E8A1EC7A7AAAFA191DFCD24732991CCA4CE081485ECE";
    attribute INIT_2D of inst : label is "77D56D2976C5E0938B90AD1A09431ECB6536CC49BE39D8F5256386BCC5A9E247";
    attribute INIT_2E of inst : label is "0818F9392AA66A28F8D7A4EAD2D79AB766BF8DCB8930E52AF524A6C8525F66A2";
    attribute INIT_2F of inst : label is "6E6A2AF780B4A598A7DE43B25E21A58D484645F2BCC427E7A473A7630C923351";
    attribute INIT_30 of inst : label is "6E11409BE752DACEDBA461461DD9AFA861FD2197918E8D6DB36C8A598E9F723E";
    attribute INIT_31 of inst : label is "99606AB8F4D266AA91EFBA229B66A89DA4A2084B0A872DD09CD0B39327EA1A4F";
    attribute INIT_32 of inst : label is "91EF5519775C19D7703885D1B9ED609952059E8A8B7DA1E1FDE5F52564BBDC48";
    attribute INIT_33 of inst : label is "A61D92AFCB3B3E321658EFEF8B8BBA5211DFB68AEE192B1B861D119A91D2A165";
    attribute INIT_34 of inst : label is "5E58AC762D123985C5A904DD7599ABBBA891199744A6DED1D57A869186BED577";
    attribute INIT_35 of inst : label is "7469691172ED21BBD62BBE26A572E16F8B84A524A95DB84662AB08F316582E1E";
    attribute INIT_36 of inst : label is "8B8456D6D7FF115B885F5B4A4757654460647347769D84AB6A91A564A4108291";
    attribute INIT_37 of inst : label is "7485871E346858291D219E2D51AB44745692D6CBA25B898A6DACBA623EE1F125";
    attribute INIT_38 of inst : label is "B528F5814AC8A213896585A2C7C787965B1E7920ADD44106791CB6B75D1769D7";
    attribute INIT_39 of inst : label is "6DE4418A271A79EC6CA7828116CD3B3A3478176DE8B1BBC49618792D6D25B6A5";
    attribute INIT_3A of inst : label is "C7521B1EBC7C7E32F2F8931256C6185F889961F8925C797D7D25B1E78086DA7C";
    attribute INIT_3B of inst : label is "C7D6C3186D248380971E7B44386D646C29E92D20B2B7434282CE87C2087DE787";
    attribute INIT_3C of inst : label is "B5B1F39FDA010471F7D21B0F482D2160B5D207D49758BD39B484D2096171FD25";
    attribute INIT_3D of inst : label is "9707DF0628793C2034971C4D617DF4B7F3B7B3B383F2920ACE0BDB2821ACA0B0";
    attribute INIT_3E of inst : label is "8FFAFBF7EB2C6B7B39E0B1A0B7B0B4B3B0B0B6F7F387DB1F125B7C707D3D61F0";
    attribute INIT_3F of inst : label is "3C0D71F4C4C4C4C0D7C717DF025F0B5F1E438C1F6C4485F4B1868382C6F383B2";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "01B866E43A3E2523EC1C0B310028809EF48A6AE137071120080800001D510458";
    attribute INIT_01 of inst : label is "C7DB47F037FA32611C74D59BD17B1137DAABAAE3AFC2337CE1917FAA344B14B7";
    attribute INIT_02 of inst : label is "8062F85BF40A5F82D9C68064A9A4B2402CB1F4DE3799D5BADC0465327B214153";
    attribute INIT_03 of inst : label is "FBFF257D49A66E49C2C02B557BD58C8B16B140F6D672BDD282F83B8F6449D11D";
    attribute INIT_04 of inst : label is "124EAED0ED16EC01E386298FD3639D219F7E42ADDF1B203E57DF832B6328AD28";
    attribute INIT_05 of inst : label is "8302CA77CE4524E8013B0EF90C87646F72409DBA3A1B76C8D879A289C60C6EE2";
    attribute INIT_06 of inst : label is "3E211EDD12961FA6C6356EC28FECF291CA54D6B8E1AF883988E348E02DFD765B";
    attribute INIT_07 of inst : label is "8E6A88D42FB671890751E5047F44D254CD84941DA5A44A75337CD213BC0AB0BF";
    attribute INIT_08 of inst : label is "6221B56981C0DD25C9813DABF7B55475C79A80E1821217729091FF9035D69BBE";
    attribute INIT_09 of inst : label is "BC9AB4EDE0D8CB3FA316EF196887DE74127A007F5D06796363E393027F593274";
    attribute INIT_0A of inst : label is "AB4B5C99ED2EAE8314F30BC293334AFECD555F7B35E61E9AA07970CB7961E9EB";
    attribute INIT_0B of inst : label is "6AC8E720D8B3AEF4F4D0DDE7763EC1753BF2CAB12B3C8FA6F02C9DA4F0003913";
    attribute INIT_0C of inst : label is "F24E2FC71A557A79581674EA7F7BB252A5D2AD9BB0D6C0E4B0607427C841E178";
    attribute INIT_0D of inst : label is "844D79B43942AB3EDD54FB63E002A442C0FAFA234F1E8D652AA2B60D43A20B4A";
    attribute INIT_0E of inst : label is "5B144B2C5E08FDFDF4596149BD2920FCDFFCB7EC551ADCF0BA0C8F0294C4FDB0";
    attribute INIT_0F of inst : label is "446AA7F48052ED417EF6823CBD9D26BCC851F9383F407143C7F3C9EAA196AF85";
    attribute INIT_10 of inst : label is "3F11592AE85A697311344BB8E7DCDCD13CB364208863E95B3D76724B4556227A";
    attribute INIT_11 of inst : label is "6599AA9F21EF494AD25A38E6BA8884C5D88529510B10949EB95AB2A79EA51F70";
    attribute INIT_12 of inst : label is "99A38EBA6A2BB7A21058377E9EDD75929A430AD824074928A94669481E47FF48";
    attribute INIT_13 of inst : label is "80D9D4FDCC7AD8F5AE412B0CFAD6188693174C6032918A98EA4C76E1E5B17D37";
    attribute INIT_14 of inst : label is "97BF5301949C0770FB132F0B6417EB9B95775B7EAD9C45EB2774B827D1EAD746";
    attribute INIT_15 of inst : label is "290D154033B487110CCF79EAE3EF8BDD39C07A7E0BF83E5C47FEECA0C0BDDDC0";
    attribute INIT_16 of inst : label is "5B5E8872DEFB3A5D21CDD7708D3E2C0DD7704E5184A20FFA2C3056D4C7FBDF01";
    attribute INIT_17 of inst : label is "4CFB862898A6C3F3DE7C533CF4A7AFD679CC39186E19687035A2F29749D87039";
    attribute INIT_18 of inst : label is "66587DE0F19A86203C2597B55A481A71FDF30C3492C1E71E7933F4C341A83C93";
    attribute INIT_19 of inst : label is "29A69186687D296D6A60E9897A3F59A4A290E65FA1B92C969245142687A5A49E";
    attribute INIT_1A of inst : label is "965D55152A2AA4466679AD66679E7A7B6DB60975586A87814814665785496649";
    attribute INIT_1B of inst : label is "4A5665D18484861915ED5A9A549255E5A1E12D5A97AEBA88612B98A61B61ED66";
    attribute INIT_1C of inst : label is "A2A6AA955B47786E647B86AE861D5545E7AA5D144A9524AEABAD2D2D145265A8";
    attribute INIT_1D of inst : label is "B51B4B696AADE1EBB787AE8B4AE1EBB452D1D518AAE18A2BAAE87B4446D62BAE";
    attribute INIT_1E of inst : label is "4921FB91D257186D22BADEB9E1A4B546D21E1D1E2E4878786DB6AAA9692DE1A5";
    attribute INIT_1F of inst : label is "E4B7B4B78791DBAB792D21E1A4B5B492C61F4B5B7EB792BB4B7879E1E0F4F492";
    attribute INIT_20 of inst : label is "792D64B4B182D21E5F486DED2DE1E1E1E78796D61B0B48692C61A1E492086DAD";
    attribute INIT_21 of inst : label is "6C2DB7861B1A082C2CE7B086DB1F79E0B686C2D2D24B7DFD2DE1F1FBB783C3DF";
    attribute INIT_22 of inst : label is "83C7C49F1E02187C3C2CF7C0931F12493D21F4F48487DF7C27B4B4C4921B787C";
    attribute INIT_23 of inst : label is "F7DF7820B7C092087C3C3DE4B082C2C21B780821B7B38782C2824B183DF4B3B7";
    attribute INIT_24 of inst : label is "2C2CE0E0F1FDF1E0F0F7C31FDE0821F1EDF020F087D3024C71F1F7DF0F0860F0";
    attribute INIT_25 of inst : label is "3DF48303030F0F7D3037C30F0C30C3C3CF0F0F7C083C2C2CF0B0FCF38E0F3DEC";
    attribute INIT_26 of inst : label is "3F08FCF7C23C3C3CF082CFCF0C2CF0F0F7B083C30C30F0F0F3C3020B0F0F4C30";
    attribute INIT_27 of inst : label is "0F3F083C30C30F7C3C7DF030D3037F0830F7C083C3C3C3C3DF0831C7CF3F3C7F";
    attribute INIT_28 of inst : label is "0F7C3C083C30C3CF3C3CF0B3C3C2CF7F0F0C20F3CFC3DF0F7F083CF3C20F0B0F";
    attribute INIT_29 of inst : label is "FCF7F38FCF7F0F0C30F0C3CF0C30F0C303DF0F0F4C3C7C3C0C3C31F0C3C3CF0F";
    attribute INIT_2A of inst : label is "F09303C3C30F030F1C3C3C3C3C30F0C0DFC3CFCF383C3DF3C3C3C3CF7C0C3F3D";
    attribute INIT_2B of inst : label is "C20F0C2C3CF3C20C3DFCF3C3C20FCF0C3C7C30C3C3F3C0C31F0F0F0F7C30F0F7";
    attribute INIT_2C of inst : label is "B1F7C7C3C30C3DF0C3C3C3C3CF0F0F0F3C30C3CF0C30F0F0C3C3DFC30C3DFCF3";
    attribute INIT_2D of inst : label is "C2C30F0F0FDFC30F3F3C383C3C30FCF3F0F083C3F3F083CF0F0F0C2C3C3C3C30";
    attribute INIT_2E of inst : label is "30C3CF0F0F0F0F7C3C0F0C3CF0F0F0F0F7F3C083DF03C303C3030F0C0C3CF0F7";
    attribute INIT_2F of inst : label is "0F0F0F3F0C3C3C3C3CFC30F0F3C3C3C3C3C3C3CFCFC30F3F3C3F3F3C3C30F0F0";
    attribute INIT_30 of inst : label is "F3C30C3F3F0CFCFCF3C30F0C3C3C3CF0C3CF030F0C3C3C30F0F0C0C3C3C3C30F";
    attribute INIT_31 of inst : label is "C0C30F3C3C0F0F3CF0F3CF030F0F3C3C3DF030C3C3C3CFC3CFC33F0F0F3C3C3C";
    attribute INIT_32 of inst : label is "F0F3C30F3F083CF3F0F3C3C3CFCF0C3C30C3C3C3C3CFC3C3CFC3C3030C3CF0C0";
    attribute INIT_33 of inst : label is "3C3C30F3C30F0F03030C3CF3C3C3CF0C30F3F0C3CF030F0F0C3C303CF0F0F0F0";
    attribute INIT_34 of inst : label is "0F0C3C3C3C30F3C3C3CF0CFCF3CF3F3CF0C30F0F0C3CFCF0F0F3C3C3C3CFC30F";
    attribute INIT_35 of inst : label is "3C3C3C30F0FC30F3C30F3C30F0F0F033C3C0C30C3C3C3C0C30F300C3030C0F0F";
    attribute INIT_36 of inst : label is "C3C0C3C3C3CF030F0C0F0F0F0F0F3C30F0F0F3C3F3CF0C3F3CF0F0F0F0C3C3C3";
    attribute INIT_37 of inst : label is "F0C3C3CF3C3C3C3C3C30FC3C30F3C0F0C3C3C3C3C30F0C0C3C3C3C303CF0F030";
    attribute INIT_38 of inst : label is "F030F0C0C3C0C3030C30C0C3C3C3C3C30F0F3C30FCF0C30F3C3CF3F3CF0F3CF3";
    attribute INIT_39 of inst : label is "3CF0C3CF3F0F3CFC3CF3C3C30FCF3F3F3C3C0F3CF0F0F3C0C30C3C3C3C30F0F0";
    attribute INIT_3A of inst : label is "C3C30F0F3C3C3C30F0F0C30303C30C0F0C0C30F0C30C3C3C3C30F0F3C0C3CF3C";
    attribute INIT_3B of inst : label is "C3C3C30C3C30C3C0C30F3F0C3C3C3C3C3CFC3C30F3F3C3C3C3CFC3C30C3CF3C3";
    attribute INIT_3C of inst : label is "F3F3F3CFCF030C30F3C30F0F0C3C3030F0C303C0C30C3C30F0C0C30C3030FC30";
    attribute INIT_3D of inst : label is "C303CF030C3C3C3030C30C0C303CF0F3F3F3F3F3C3F3C30FCF0FCF3C30FCF0F0";
    attribute INIT_3E of inst : label is "CFFFFFFFFF3C3F3F3CF0F0F0F3F0F0F3F0F0F3F3F3C3CF0F030F3C303C3C30F0";
    attribute INIT_3F of inst : label is "3C0C30F0C0C0C0C0C3C303CF030F0F0F0F030C0F3C00C0F0F0C3C3C3C3F3C3F3";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "5B455475A4B7861B6AE492C6D61B1F79E1F0F0F03308BA0009090001BA110B01";
    attribute INIT_01 of inst : label is "ED57B91211A1851E84A96EA462D1B95451565451A1491B9EABAEB7455EE1EB91";
    attribute INIT_02 of inst : label is "5BBAAA17762AE9546AEB62B55EA5455BAE46927569EB4AD744A2A5854515BB95";
    attribute INIT_03 of inst : label is "D445455146446A86A26E145515EAEA552AD9197B55191EB9E114A926AE546E85";
    attribute INIT_04 of inst : label is "EBAAB5E85EB97AEBD6BAA85AADB914A857A46EB547A05675276D55291AA16BAA";
    attribute INIT_05 of inst : label is "A854AAAAA94A850AEA4685DBAE45B6F5DEBE514497ADBA5156E97AE549249E7A";
    attribute INIT_06 of inst : label is "0518A4264867E76E5294AA71457A51491BD91498519B6EB646E94AABAAAA5E97";
    attribute INIT_07 of inst : label is "A517E454E0297ABA152A3A8615F9A1685155BA914685551A45146EAAD68519DA";
    attribute INIT_08 of inst : label is "BAB91682AE4946EA152BA517D429A1951BA5FAD85BE46AAB6A7E242A452AAA90";
    attribute INIT_09 of inst : label is "E5494660527E129769F57682946E6D9EA7D685B952A7D46AAB546EA15829AE45";
    attribute INIT_0A of inst : label is "1AE4667D6457A45BD6E9B991A0D9857682AE5F597D2F660A4057A9F5AAB97D65";
    attribute INIT_0B of inst : label is "825BA45BA51A60651BA52606B6960D6B975C1ACD9B84A5825A775F5A3E6F916F";
    attribute INIT_0C of inst : label is "5F90D585919B97D685551A60911AA82AA82AA43594A6535A0A52AE84BDAE9196";
    attribute INIT_0D of inst : label is "61867A5F97EB679E7ABAD45452B146BABAD8119F661436DA825452A0A814DDBD";
    attribute INIT_0E of inst : label is "A0A866DE45245E76B6452A145E82A158275E7982B927D4525EA15159F67E76D8";
    attribute INIT_0F of inst : label is "4920850A86482619109E49279E45679F7AEB9EA19D4EABAE79E9E8149EBD46AE";
    attribute INIT_10 of inst : label is "90921857986DE49F61F649B609B605249B79F64867D82D9EA9149F67AE48679E";
    attribute INIT_11 of inst : label is "B79279E086DA49F60879F609E7921921B4924861F7DF486D821B6DE4B609209F";
    attribute INIT_12 of inst : label is "7927920B7920B7861F4926C2D82DE4879F7C36DB4936D21B7921821860869B61";
    attribute INIT_13 of inst : label is "DF083DE083C2082DE087DB79E6DE487D86DF7921F6D21B79209F6DE49F61824B";
    attribute INIT_14 of inst : label is "DE0B7C7DF7D87C21E0F7C21821F782DE7DE7DE08209F7DE0F6092D279F0820F7";
    attribute INIT_15 of inst : label is "C3DF7DF1F6C3DF7C7D820820B782DE092DF7C20B482D2083D23839F7DF082087";
    attribute INIT_16 of inst : label is "7CF3DF0F082C20F0F7D83C21F0F3C3183C21F0F7DF0F48E0F0C37C3DF0820837";
    attribute INIT_17 of inst : label is "3DE0F0C3C30F0F3CF3CF0C2083C20B3C209F0F7DF3C3C3C30F0F3C3C3083C30F";
    attribute INIT_18 of inst : label is "F0F0CFC33C3C30C30F0F0F3C3C30C3C3CF3C30C30F0C3C33CF7F3DF0C7C30F0C";
    attribute INIT_19 of inst : label is "0F0F0C30F0CF0F0F0F0C3C30F0F3C3C30F0C3C3CF7CF0F0F0C30C30F0F3C3C3C";
    attribute INIT_1A of inst : label is "0C3C30C30F0F3C30F0F3CF0F0F3CF3F3CF3C30F0C30F0F0C30C30F0F0C30F0C3";
    attribute INIT_1B of inst : label is "C3C3C3C30C0C0C30C3CF0F0F0C30C3C3C3C30F0F0F3CF3C0C30F3C3C33C3CF0F";
    attribute INIT_1C of inst : label is "F0F0F3C30F0F3C3CF0F3C3CF0C3C30C3CF3C3C30C3C30C3CF3CF0F0F0C30F0F0";
    attribute INIT_1D of inst : label is "F30F0F3C3CFCF0F3F3C3CF0F0CF0F3F0C3C3C30C3CF0C30F3CF0F3C0C3C30F3C";
    attribute INIT_1E of inst : label is "0C30F3C3C30F0C3C30F3CF3CF0F0F0C3C30F0F0F0F0C3C3C3CF3CF3C3C3CF0F0";
    attribute INIT_1F of inst : label is "F0F3F0F3C3C3CF3F3C3C30F0F0F0F0C3C30F0F0F3CF3C33F0F3C3CF0F0F0F0C3";
    attribute INIT_20 of inst : label is "3C3C30F0F0C3C30F0F0C3CFC3CF0F0F0F3C3C3C30F0F0C3C3C30F0F0C30C3CFC";
    attribute INIT_21 of inst : label is "3C3CF3C30F0F0C3C3CF3F0C3CF0F3CF0F3C3C3C3C30F3CFC3CF0F0F3F3C3C3CF";
    attribute INIT_22 of inst : label is "C3C3C0CF0F030C3C3C3CF3C0C30F030C3C30F0F0C0C3CF3C33F0F0C0C30F3C3C";
    attribute INIT_23 of inst : label is "F3CF3C30F3C0C30C3C3C3CF0F0C3C3C30F3C0C30F3F3C3C3C3C30F0C3CF0F3F3";
    attribute INIT_24 of inst : label is "3C3CF0F0F0FCF0F0F0F3C30FCF0C30F0FCF030F0C3C3030C30F0F3CF0F0C30F0";
    attribute INIT_25 of inst : label is "3CF0C303030F0F3C3033C30F0C30C3C3CF0F0F3C0C3C3C3CF0F0FCF3CF0F3CFC";
    attribute INIT_26 of inst : label is "3F0CFCF3C33C3C3CF0C3CFCF0C3CF0F0F3F0C3C30C30F0F0F3C3030F0F0F0C30";
    attribute INIT_27 of inst : label is "0F3F0C3C30C30F3C3C3CF030C3033F0C30F3C0C3C3C3C3C3CF0C30C3CF3F3C3F";
    attribute INIT_28 of inst : label is "0F3C3C0C3C30C3CF3C3CF0F3C3C3CF3F0F0C30F3CFC3CF0F3F0C3CF3C30F0F0F";
    attribute INIT_29 of inst : label is "FCF3F3CFCF3F0F0C30F0C3CF0C30F0C303CF0F0F0C3C3C3C0C3C30F0C3C3CF0F";
    attribute INIT_2A of inst : label is "F0C303C3C30F030F0C3C3C3C3C30F0C0CFC3CFCF3C3C3CF3C3C3C3CF3C0C3F3C";
    attribute INIT_2B of inst : label is "C30F0C3C3CF3C30C3CFCF3C3C30FCF0C3C3C30C3C3F3C0C30F0F0F0F3C30F0F3";
    attribute INIT_2C of inst : label is "F0F3C3C3C30C3CF0C3C3C3C3CF0F0F0F3C30C3CF0C30F0F0C3C3CFC30C3CFCF3";
    attribute INIT_2D of inst : label is "C3C30F0F0FCFC30F3F3C3C3C3C30FCF3F0F0C3C3F3F0C3CF0F0F0C3C3C3C3C30";
    attribute INIT_2E of inst : label is "30C3CF0F0F0F0F3C3C0F0C3CF0F0F0F0F3F3C0C3CF03C303C3030F0C0C3CF0F3";
    attribute INIT_2F of inst : label is "0F0F0F3F0C3C3C3C3CFC30F0F3C3C3C3C3C3C3CFCFC30F3F3C3F3F3C3C30F0F0";
    attribute INIT_30 of inst : label is "F3C30C3F3F0CFCFCF3C30F0C3C3C3CF0C3CF030F0C3C3C30F0F0C0C3C3C3C30F";
    attribute INIT_31 of inst : label is "C0C30F3C3C0F0F3CF0F3CF030F0F3C3C3CF030C3C3C3CFC3CFC33F0F0F3C3C3C";
    attribute INIT_32 of inst : label is "F0F3C30F3F0C3CF3F0F3C3C3CFCF0C3C30C3C3C3C3CFC3C3CFC3C3030C3CF0C0";
    attribute INIT_33 of inst : label is "3C3C30F3C30F0F03030C3CF3C3C3CF0C30F3F0C3CF030F0F0C3C303CF0F0F0F0";
    attribute INIT_34 of inst : label is "0F0C3C3C3C30F3C3C3CF0CFCF3CF3F3CF0C30F0F0C3CFCF0F0F3C3C3C3CFC30F";
    attribute INIT_35 of inst : label is "3C3C3C30F0FC30F3C30F3C30F0F0F033C3C0C30C3C3C3C0C30F300C3030C0F0F";
    attribute INIT_36 of inst : label is "C3C0C3C3C3CF030F0C0F0F0F0F0F3C30F0F0F3C3F3CF0C3F3CF0F0F0F0C3C3C3";
    attribute INIT_37 of inst : label is "F0C3C3CF3C3C3C3C3C30FC3C30F3C0F0C3C3C3C3C30F0C0C3C3C3C303CF0F030";
    attribute INIT_38 of inst : label is "F030F0C0C3C0C3030C30C0C3C3C3C3C30F0F3C30FCF0C30F3C3CF3F3CF0F3CF3";
    attribute INIT_39 of inst : label is "3CF0C3CF3F0F3CFC3CF3C3C30FCF3F3F3C3C0F3CF0F0F3C0C30C3C3C3C30F0F0";
    attribute INIT_3A of inst : label is "C3C30F0F3C3C3C30F0F0C30303C30C0F0C0C30F0C30C3C3C3C30F0F3C0C3CF3C";
    attribute INIT_3B of inst : label is "C3C3C30C3C30C3C0C30F3F0C3C3C3C3C3CFC3C30F3F3C3C3C3CFC3C30C3CF3C3";
    attribute INIT_3C of inst : label is "F3F3F3CFCF030C30F3C30F0F0C3C3030F0C303C0C30C3C30F0C0C30C3030FC30";
    attribute INIT_3D of inst : label is "C303CF030C3C3C3030C30C0C303CF0F3F3F3F3F3C3F3C30FCF0FCF3C30FCF0F0";
    attribute INIT_3E of inst : label is "CFFFFFFFFF3C3F3F3CF0F0F0F3F0F0F3F0F0F3F3F3C3CF0F030F3C303C3C30F0";
    attribute INIT_3F of inst : label is "3C0C30F0C0C0C0C0C3C303CF030F0F0F0F030C0F3C00C0F0F0C3C3C3C3F3C3F3";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "A5A69A5A5A5969A5965A696969A5A5965A5A5A5A990255000000000015550255";
    attribute INIT_01 of inst : label is "65A5969A9A5A69A5A696965A6969969A69A5A69A5A69A596596595A6965A5969";
    attribute INIT_02 of inst : label is "A59659A5969965A696596996965A69A59669699696596965A69A5A69A69A5969";
    attribute INIT_03 of inst : label is "5A69A69A69A6966969969A69A65965A699669A5969A6965969A6969965A69669";
    attribute INIT_04 of inst : label is "65965966965996596659669965969A6699669659A59A69969965A699A59A6596";
    attribute INIT_05 of inst : label is "669A659659A669A659A6696596699659659669A699659669A659965A69A69659";
    attribute INIT_06 of inst : label is "A69A6699A6996596699A659A699669A699669A669A659659A659A65965966599";
    attribute INIT_07 of inst : label is "6699669A66999659A6999669A6599A669A699669A669A699A69A65996669A659";
    attribute INIT_08 of inst : label is "9659A6699669A659A699669966999A66996659669966996599966699A699659A";
    attribute INIT_09 of inst : label is "59A6699A69966999665996699A6596659966699669996699659A659A66999669";
    attribute INIT_0A of inst : label is "9966999666996699665996699A66699669966599966599A66A99665996599666";
    attribute INIT_0B of inst : label is "6999669966999A66996699A65999A66599669966659A66699996659996659A65";
    attribute INIT_0C of inst : label is "659A66699A65996669A6999A66996699669966999A666999A669966996659A66";
    attribute INIT_0D of inst : label is "9A699665996599659659669A699A699659669A6599A69966699A699A669A6596";
    attribute INIT_0E of inst : label is "9A669965A69A659659A699A696699A66996596699699669A659A69A659965966";
    attribute INIT_0F of inst : label is "A69A69A669A699A69A65A69965A699659659659A65A659659659669A65966965";
    attribute INIT_10 of inst : label is "9A69A69966965A659A59A659A659A69A659659A699669665969A659965A69965";
    attribute INIT_11 of inst : label is "5969965A6965A659A69659A65969A69A5A69A69A5965A69669A5965A59A69A65";
    attribute INIT_12 of inst : label is "969969A5969A5969A5A6996966965A6965969965A69969A5969A69A69A69659A";
    attribute INIT_13 of inst : label is "65A6965A6969A6965A6965965965A6966965969A5969A5969A65965A659A69A5";
    attribute INIT_14 of inst : label is "65A596965966969A5A5969A69A596965965965A69A65965A59A6969965A69A59";
    attribute INIT_15 of inst : label is "6965965A596965969669A69A596965A6965969A5A6969A696996965965A69A69";
    attribute INIT_16 of inst : label is "965965A5A6969A5A5966969A5A5969A6969A5A5965A5A65A5A6996965A69A699";
    attribute INIT_17 of inst : label is "965A5A6969A5A5965965A69A6969A5969A65A59659696969A5A596969A6969A5";
    attribute INIT_18 of inst : label is "5A5A656996969A69A5A5A596969A696965969A69A5A696996595965A6969A5A6";
    attribute INIT_19 of inst : label is "A5A5A69A5A65A5A5A5A6969A5A596969A5A696965965A5A5A69A69A5A5969696";
    attribute INIT_1A of inst : label is "A6969A69A5A5969A5A5965A5A596595965969A5A69A5A5A69A69A5A5A69A5A69";
    attribute INIT_1B of inst : label is "69696969A6A6A69A6965A5A5A69A69696969A5A5A596596A69A59696996965A5";
    attribute INIT_1C of inst : label is "5A5A5969A5A596965A596965A6969A696596969A6969A6965965A5A5A69A5A5A";
    attribute INIT_1D of inst : label is "59A5A59696565A59596965A5A65A595A696969A6965A69A5965A596A6969A596";
    attribute INIT_1E of inst : label is "A69A596969A5A6969A5965965A5A5A6969A5A5A5A5A696969659659696965A5A";
    attribute INIT_1F of inst : label is "5A595A596969659596969A5A5A5A5A6969A5A5A596596995A596965A5A5A5A69";
    attribute INIT_20 of inst : label is "96969A5A5A6969A5A5A69656965A5A5A59696969A5A5A696969A5A5A69A69656";
    attribute INIT_21 of inst : label is "96965969A5A5A69696595A6965A5965A5969696969A59656965A5A5959696965";
    attribute INIT_22 of inst : label is "69696A65A5A9A6969696596A69A5A9A6969A5A5A6A696596995A5A6A69A59696";
    attribute INIT_23 of inst : label is "5965969A596A69A69696965A5A696969A596A69A595969696969A5A6965A5959";
    attribute INIT_24 of inst : label is "96965A5A5A565A5A5A5969A565A69A5A565A9A5A6969A9A69A5A5965A5A69A5A";
    attribute INIT_25 of inst : label is "965A69A9A9A5A5969A9969A5A69A696965A5A596A69696965A5A565965A59656";
    attribute INIT_26 of inst : label is "95A65659699696965A696565A6965A5A595A6969A69A5A5A5969A9A5A5A5A69A";
    attribute INIT_27 of inst : label is "A595A6969A69A59696965A9A69A995A69A596A696969696965A69A6965959695";
    attribute INIT_28 of inst : label is "A59696A6969A696596965A5969696595A5A69A59656965A595A6965969A5A5A5";
    attribute INIT_29 of inst : label is "565959656595A5A69A5A6965A69A5A69A965A5A5A6969696A6969A5A696965A5";
    attribute INIT_2A of inst : label is "5A69A96969A5A9A5A6969696969A5A6A65696565969696596969696596A69596";
    attribute INIT_2B of inst : label is "69A5A696965969A69656596969A565A696969A6969596A69A5A5A5A5969A5A59";
    attribute INIT_2C of inst : label is "5A59696969A6965A6969696965A5A5A5969A6965A69A5A5A69696569A6965659";
    attribute INIT_2D of inst : label is "6969A5A5A56569A595969696969A56595A5A6969595A6965A5A5A6969696969A";
    attribute INIT_2E of inst : label is "9A6965A5A5A5A59696A5A6965A5A5A5A59596A6965A969A969A9A5A6A6965A59";
    attribute INIT_2F of inst : label is "A5A5A595A696969696569A5A59696969696969656569A59596959596969A5A5A";
    attribute INIT_30 of inst : label is "5969A69595A656565969A5A69696965A6965A9A5A696969A5A5A6A69696969A5";
    attribute INIT_31 of inst : label is "6A69A59696A5A5965A5965A9A5A59696965A9A6969696569656995A5A5969696";
    attribute INIT_32 of inst : label is "5A5969A595A696595A5969696565A6969A69696969656969656969A9A6965A6A";
    attribute INIT_33 of inst : label is "96969A5969A5A5A9A9A69659696965A69A595A6965A9A5A5A6969A965A5A5A5A";
    attribute INIT_34 of inst : label is "A5A69696969A59696965A656596595965A69A5A5A696565A5A596969696569A5";
    attribute INIT_35 of inst : label is "9696969A5A569A5969A5969A5A5A5A99696A69A6969696A69A59AA69A9A6A5A5";
    attribute INIT_36 of inst : label is "696A69696965A9A5A6A5A5A5A5A5969A5A5A59695965A695965A5A5A5A696969";
    attribute INIT_37 of inst : label is "5A69696596969696969A56969A596A5A6969696969A5A6A69696969A965A5A9A";
    attribute INIT_38 of inst : label is "5A9A5A6A696A69A9A69A6A6969696969A5A5969A565A69A59696595965A59659";
    attribute INIT_39 of inst : label is "965A696595A5965696596969A56595959696A5965A5A596A69A69696969A5A5A";
    attribute INIT_3A of inst : label is "6969A5A59696969A5A5A69A9A969A6A5A6A69A5A69A69696969A5A596A696596";
    attribute INIT_3B of inst : label is "696969A6969A696A69A595A6969696969656969A5959696969656969A6965969";
    attribute INIT_3C of inst : label is "5959596565A9A69A5969A5A5A6969A9A5A69A96A69A6969A5A6A69A69A9A569A";
    attribute INIT_3D of inst : label is "69A965A9A696969A9A69A6A69A965A5959595959695969A565A565969A565A5A";
    attribute INIT_3E of inst : label is "6555555555969595965A5A5A595A5A595A5A5959596965A5A9A5969A96969A5A";
    attribute INIT_3F of inst : label is "96A69A5A6A6A6A6A6969A965A9A5A5A5A5A9A6A596AA6A5A5A69696969596959";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
