-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FA66D24D0DD03021E6799E79A0864247FFFB315A69EE80EFFFF1FEB3E7FFFF6D";
    attribute INIT_01 of inst : label is "99A559CC99DF17C5F8DB34A6404D468BD61234FC1382F7578002CAE1AB71F7D7";
    attribute INIT_02 of inst : label is "1743F1EBB88F9C6C204C433067763840551C4B30AA8802BD856FBE93D7A9EBB4";
    attribute INIT_03 of inst : label is "11A20AA1CC2D7D7A4AAE42B0F07A7871E02EEAFD8E77CC243D3BE060C465A1DF";
    attribute INIT_04 of inst : label is "40148A2890120B4D658448535565E3CF0E34000AC228452800044449810A1341";
    attribute INIT_05 of inst : label is "DB0A616913140519143814AC0B6A1C738EF12A854D4C844461702B60938B4A8B";
    attribute INIT_06 of inst : label is "DB501003FD57F63F6AF77D4008A28BFEBEA37B725AE313C2C6F25DF1217BA4D4";
    attribute INIT_07 of inst : label is "E2044DFF16B0CE2FA25A098131596592A825925AB96A4CA0A14537392160DE79";
    attribute INIT_08 of inst : label is "DFBD224E9A9BB04920036E0B92ADBC8AB77F0935C031D11F0988AC0B5D8382C0";
    attribute INIT_09 of inst : label is "E3214CC0543709044C9BA7F2E9FC9DDA7FC0FA41810F52EF84804C0EC4A0144C";
    attribute INIT_0A of inst : label is "999BFB6085CC1C4F6F347FBDB480246A16ACA339773B2CDD0ABEC4158850A028";
    attribute INIT_0B of inst : label is "21E2605020107F5ADAD2AE974BA4E89800B45C12E69346DB2F3210D64F00A85F";
    attribute INIT_0C of inst : label is "1B1D5C961304E92F92F96F962CACBE26BEBB3B39ACABDBD24FE3470E0C00C360";
    attribute INIT_0D of inst : label is "2236FA046D96CD75D2184C6A1BD24EABDB2DF7A0F45DE9ABC8672938A715A706";
    attribute INIT_0E of inst : label is "4A1A1CF8A74E026F3B3554D9D488E6EC0C11AE90D4A0D3CEAC5A63C7A6134931";
    attribute INIT_0F of inst : label is "EA602A8003B40AA000ED0640440549D39F375E3BF67CFBAAE66033BC3BB9CFE8";
    attribute INIT_10 of inst : label is "80155D41614C2CE671B75C67DD2B7EEB0E2CC4C5E84B3B26FC622200206397D9";
    attribute INIT_11 of inst : label is "C63E64E4727194669055241432EAA82404009002184A13FFAB241F27C1227BF3";
    attribute INIT_12 of inst : label is "067D18B75E0CD1C899782A4888AD34A405E00000008020080204C18616CA8E02";
    attribute INIT_13 of inst : label is "393137F610935206CA23210EE6F60A64FA42103999E7891E02C6FE81330A54CC";
    attribute INIT_14 of inst : label is "595F8C0A059603E109249A8B220411170100410D93411156490498361424261F";
    attribute INIT_15 of inst : label is "51150DC0822B4AC8AC94885B23F52AD4203466BDA730B399FBAD09CB1B6CC7EC";
    attribute INIT_16 of inst : label is "6659043B21A3A30E8993370A6F734A8A49626E3062951648E16078B4B1301772";
    attribute INIT_17 of inst : label is "02081E1E7DF91E0656B4B6BE71E2C92083D8230C0B096F5993841882CF0A620A";
    attribute INIT_18 of inst : label is "2184F73CF164F2D301BAE458E290231C192625F29EB96B1C9D855BC9080AC896";
    attribute INIT_19 of inst : label is "028EB24D671692C080FBE00A05FBACF8EC40206B5F820180002A200419B8CB04";
    attribute INIT_1A of inst : label is "400010003B3ECFF700000000001000804E60659675EFFAFE4C8BEFEBE7D84FAC";
    attribute INIT_1B of inst : label is "00000200FB58DFF6000000002050112010001000D53FDF370000000004E60225";
    attribute INIT_1C of inst : label is "3C0CB0844D4405C08C209424924856B41584DA724861FC8D6A81771C624076EB";
    attribute INIT_1D of inst : label is "F55FF505588180186C7878FADA908172EE1570313D051ADCE1E7C7A1D015E20C";
    attribute INIT_1E of inst : label is "B1D1D2A8DA5F90011033198A0C21C8C4D8130ACDD65F592F0646224308510510";
    attribute INIT_1F of inst : label is "F3F0DDFEFBFEF3E64000180400000000F5CAE7D635BE057B0000000000000000";
    attribute INIT_20 of inst : label is "229D4EBEB712660301C0EB7539CCB239B88E33331C5011114469B9B336E62608";
    attribute INIT_21 of inst : label is "FEBD9E72782733F9AB295465BCD56C95D4A66A3BBBB8D4DE6D64DA9D0D524BB5";
    attribute INIT_22 of inst : label is "83001020831D90B38EF7139A931F0567CDD78EFD9FC987B2EC0277AD91F5098F";
    attribute INIT_23 of inst : label is "40100C022008A80AC82082CE80028688A0200028031145101150571005445575";
    attribute INIT_24 of inst : label is "90402A362100448005E2F07820600F04D00480E2054015408001044640D05540";
    attribute INIT_25 of inst : label is "9C6680D0F3939F2300000000000800012000315A7FDFEFEA0000000018001D22";
    attribute INIT_26 of inst : label is "30800108D3FC6F8F000000000010400312A851417EFF5FB60000000800040800";
    attribute INIT_27 of inst : label is "274470C0A84A42E22522E9F1E7C71E1EE736360304159098578410AA4144F3DF";
    attribute INIT_28 of inst : label is "F0B971E7CF2B0CCAE58E5AC729402083ECA384B28AEBCCCC2A0B6A884849CBAF";
    attribute INIT_29 of inst : label is "44AC324B08AD22B129EC84444829F734D61401382A048903606010842B171C38";
    attribute INIT_2A of inst : label is "9B960040B0A22008B66F0565C1814000938365C918902249050801130D8946B1";
    attribute INIT_2B of inst : label is "E3F736C17E2E927E1C6987618181CCCB7CBF50502C0D215350B1525C0C32AC6F";
    attribute INIT_2C of inst : label is "7148E98D999121E001151896394396FB5CEB3AC833732D4E4CE49B62FD7FF9F1";
    attribute INIT_2D of inst : label is "6B65D08CA91584417A08DF362C88AB2C455960C59BB5128840178A20AD231364";
    attribute INIT_2E of inst : label is "B9EEFFF77E7F66D7AA67A5B8175CF1F4313534202BFD5E5B88000F0000B4A54A";
    attribute INIT_2F of inst : label is "F1F0DDDEFBEEF3E60000180400000000E54AE7D614B6256AF668EE1EF58033F3";
    attribute INIT_30 of inst : label is "C010DAB12DAB6491CBBEFA98E7EC0A69F329D169C559719D81059F3C0460BA49";
    attribute INIT_31 of inst : label is "2000002100000010401EBF7DFE8051F776F2999015BB9B5F312C8BB6ADD9E518";
    attribute INIT_32 of inst : label is "2000010000000000FFFFFFFF0648120D4240040000000000EFFFFFFF00420088";
    attribute INIT_33 of inst : label is "2400080000000000FFFDEBFF182804030800200200000000FDFB7FBF00003243";
    attribute INIT_34 of inst : label is "A06090CAF7EFB2DE000000000080000311076840B56E7FFF0000000000100000";
    attribute INIT_35 of inst : label is "1C6EC0D0F79B9F2700000001000800010000315B7FFFEFEA0000000028000000";
    attribute INIT_36 of inst : label is "30800108D3FC6F8F000000000010400312A851417EFF5FB60000000800040800";
    attribute INIT_37 of inst : label is "F0808D23CDD3FFF3000000000000080240261008BF2C37B30000000084012000";
    attribute INIT_38 of inst : label is "20020000F59F75F8100000000012014082004200DD8B7EFC0000000000800000";
    attribute INIT_39 of inst : label is "10600180FBF6FED7000000000400014000900200FD74AF66000000002488030B";
    attribute INIT_3A of inst : label is "40001000383EC7F7000000000010008040400100EB11CB5E000000000800C002";
    attribute INIT_3B of inst : label is "00000200DB58DFB4000000002054110810001000C51EDF33000000000426022D";
    attribute INIT_3C of inst : label is "CBEFE68A77DBEDB80000000200000000959BF4CA1B1928170000001200400000";
    attribute INIT_3D of inst : label is "DDA4B31AFA1A93270000000C000000006BF6AD6FF6FEC0FC0000001000000000";
    attribute INIT_3E of inst : label is "B0D110A8DA5F9AAB04410000100000001743D6A6B4DB86688000200001000400";
    attribute INIT_3F of inst : label is "F1F0DDDEFBEEF3E60000180400000000F54AE7D615BE056A0000000400000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "06092C92F478B8A8601A060012A08754800087C42051CA0000E6EBD6E0EFFF34";
    attribute INIT_01 of inst : label is "225C147ECC09304B496C49980C3D8E04C25F000F7DEFF81E0888CF63A4EC9B6C";
    attribute INIT_02 of inst : label is "D53F37919E6062F46DFD9B3266667201E01A2D725BE96618228FFEF83C9E745B";
    attribute INIT_03 of inst : label is "3CEF6920647FB5107FF0B180E06260637B722264972205B309C5CDA4462346F3";
    attribute INIT_04 of inst : label is "648FF75E3000C605BCE9C4925B1583468C71A92958F2B4E3727362705D767BE4";
    attribute INIT_05 of inst : label is "6D24A9FB886892D4B22B901E5F8CACA594B316C988C24C3365816582340581BD";
    attribute INIT_06 of inst : label is "0456595CA1F75D75DF028AA0A002BEBFEABC88BEDCFB2038916092DA4E4C0160";
    attribute INIT_07 of inst : label is "CD3D1FF9300F1072766F979268C6C630E49B3063352D2CE409A050830DE7F37D";
    attribute INIT_08 of inst : label is "BB7030865C08328212C000215ECB252204563077AD363B02251B4C91A0A9CE0F";
    attribute INIT_09 of inst : label is "19680551C6556220FD877199DC66F0994FF6E165902D42DB0736C09D06E48CC0";
    attribute INIT_0A of inst : label is "C0409EF443C807188240955DC495478A1ED1345B903C096554241C87B129FB15";
    attribute INIT_0B of inst : label is "C4748933B58632BDBFFCCCC22336454164E6FBCF844BD4AD7C31A7D040001900";
    attribute INIT_0C of inst : label is "8C5A4EE0E1DFB69965B4D945F313607968F3337E9133FBFC0B11AE1C44444780";
    attribute INIT_0D of inst : label is "C8CA339F8D5636D342692531DFA14629901133D3C108EAE47D16C0226C0667A3";
    attribute INIT_0E of inst : label is "9E9FBBED7EDC0C0FFFC2735086C99700F1A6331A606301C32A218F1CC74A370E";
    attribute INIT_0F of inst : label is "8CE0220800BC0882002F86C6EC6D69231865FBEF5C3872FF021CE38388D38713";
    attribute INIT_10 of inst : label is "2659E3E6E7DD5DFE1D066A86081480C0D0C0C80A2B344482822664220C6CBE59";
    attribute INIT_11 of inst : label is "4B363225D912D68D221424280141394E5C45192D1333E04D744F61E4C8060204";
    attribute INIT_12 of inst : label is "67AE1EE24ACEE1EBF2899476EE4DA40F170000000000000000144F5844884499";
    attribute INIT_13 of inst : label is "0B120454A3417D1EC9776F501D25794C5CC99B1C12F939233D38187717DAB6BF";
    attribute INIT_14 of inst : label is "19B7B587BD3AB6D57345A9AA468517B5DB4CDB38FD5963F4EFB2BB3D5F6EEFD2";
    attribute INIT_15 of inst : label is "AA6200A554C56FF7151F152A45F313CC4D47C222C85961FBDFB19BD826DC8764";
    attribute INIT_16 of inst : label is "78663B1E7CF55573B56BD012800AA4C53004576A85098A751287894576776122";
    attribute INIT_17 of inst : label is "235A0A147DBBE4DCA4E99BD8FE0B70D70CF33575F6F00059E1DEA93102BE84C5";
    attribute INIT_18 of inst : label is "6AD49C9442A767A9CA530CA1CFB667F88B0A8AE583CB1485F1B9E853952D9F0C";
    attribute INIT_19 of inst : label is "E56989EFD50F710E87371D6FEF1FFE8B45C8A965604996CCC4A4D64F2B5D0656";
    attribute INIT_1A of inst : label is "00000000A40201A260000023FFEDB95906A326199C1B00802C3C19180C112938";
    attribute INIT_1B of inst : label is "080000206018000004002004FFBFFCA710000000C6430831811000208DFFEFFF";
    attribute INIT_1C of inst : label is "E9AB5DE7A1CE93AD357BBDEDB780E0418A967D56DA8517C38C2C47DE6F4941D9";
    attribute INIT_1D of inst : label is "FFF55588C3488888F270E9DFBF39580AF7BCAC94D727DE0BD3870626706C0457";
    attribute INIT_1E of inst : label is "30000000200004142A554B12EA255ACFEA77CD1FC910C0C1D34F6CCC2CB64B64";
    attribute INIT_1F of inst : label is "30408002000040007ED71D457F155F020000000980000000D6E99A3C7D3FF97D";
    attribute INIT_20 of inst : label is "D70793CD2C00040000003F15800228206B0240942115400105ECA0040000EAD3";
    attribute INIT_21 of inst : label is "73C7485A7C239701808DF8F03278FAD7E9792E9FF7F8FD6F95C70B8585F2AEA9";
    attribute INIT_22 of inst : label is "0704C0000085DD3652835197675321C6197EFBD715934C24B02A147E4BF733D8";
    attribute INIT_23 of inst : label is "45511C020208208270220AD6A2228588A220288821104550511013151544456D";
    attribute INIT_24 of inst : label is "90402210310006000B64321901E003241800127C050011130886550C40B04441";
    attribute INIT_25 of inst : label is "40000000200800401A42018AADF6F57F000000006000000808C02C0050000B42";
    attribute INIT_26 of inst : label is "000000001000200000289644DF9FFFBF000000006001310001009040FFEFD5BD";
    attribute INIT_27 of inst : label is "EF51E6CB3AFC808057F0A1C1A34E9D1AEE6FEF4860843B70FFC8864908CC7B6B";
    attribute INIT_28 of inst : label is "E3C415BB7E14151F02AA8075C4BFDD7855FABF8A087AF9C97110643BDFF1EF8B";
    attribute INIT_29 of inst : label is "EC1C4411453814E294014EEFF102103765865A3B73227CC525C6D909986178F7";
    attribute INIT_2A of inst : label is "08387789742FA85A24D392810893C00030BAFA4E79F87D1CA1934837DBFBF548";
    attribute INIT_2B of inst : label is "87688FAC52C820DE41945197D7D62858022165F5351A6B66F51764CAC5545207";
    attribute INIT_2C of inst : label is "1CBC03B5155364379CA9BDF2AB0038443D5C726012346094971B6DB0BBB669C1";
    attribute INIT_2D of inst : label is "96FFDAF05F9697A58CDE7FFEDACE57B47ABD844D8BB3473EEC9CDC599C9944D6";
    attribute INIT_2E of inst : label is "4A726C1BA8F2D20060562A040FA468C5C4C1C4C0D87BBEBCA51EF2BCD94E72F7";
    attribute INIT_2F of inst : label is "3040000A000040007AD71A554F155F82002000098000000012F1709DDC02A305";
    attribute INIT_30 of inst : label is "3123DF6A559484A7A2BEE9C611C1B3496856184D0418613837DF7A704A8432CB";
    attribute INIT_31 of inst : label is "FBFFF7FF300A10A900A4FAEB1144177D5005D09B7ECA8BE25A50B45652088A8E";
    attribute INIT_32 of inst : label is "DE3FDFFB521167500104020900000000FFBEFFEF3D0004090000030C00000000";
    attribute INIT_33 of inst : label is "FBDF7FFF22024A400008050000000000FBDFFFDDB82044880200000400000000";
    attribute INIT_34 of inst : label is "000000000000000014008041FD7FFF6F800000008084104002A04007BEFB7AD5";
    attribute INIT_35 of inst : label is "40000000200800401A40018AADF6F57F000000006000000028C024005774E7F7";
    attribute INIT_36 of inst : label is "00000000100000000028964CDFDFFFBF000000006001310001009042FFEFD5BF";
    attribute INIT_37 of inst : label is "000000009080000002014000BF6E777500000000600800000102402BFEAB6FF7";
    attribute INIT_38 of inst : label is "0000000000A0000020C230607FFE0F7F00004000000800210400480066FAAF1B";
    attribute INIT_39 of inst : label is "0000000081400009208800013BEC546C000000002A80208500400001FFFF6FA6";
    attribute INIT_3A of inst : label is "00000000208201A260000023F7CD90590000000021000040040404017FFFDAFF";
    attribute INIT_3B of inst : label is "000000204018000004002004EFBEFCA710000000C2410831811000208DFBEBFD";
    attribute INIT_3C of inst : label is "00000000000000009ED74E67ED77FF3B2000300440000000EF7F0FDFF26ECE2E";
    attribute INIT_3D of inst : label is "0000080010000000B7812FED2FB191AE90001000000000004816347787FAE915";
    attribute INIT_3E of inst : label is "3000008420000000FC07B1ADB66F543880002009000000009EFF76BFEFDDF6C0";
    attribute INIT_3F of inst : label is "3040000A000040005AD71E454F155F82002000098000000086E99A147D2FB17D";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "40AB24B25440C9C80302C0B89120C3940280899A4DBDC22EFFE8E156E0EFFF1C";
    attribute INIT_01 of inst : label is "264C98649D0B02C018644B80440100C59417002E39C7F194CC9C8BA185EC3A61";
    attribute INIT_02 of inst : label is "12DE57208C618C643250FAA144440A20BA8597A014C880AA33E040290582F0D9";
    attribute INIT_03 of inst : label is "99EFCC4C26C2B1031552614A189210117171A1F4176025310B9828A62302B7C7";
    attribute INIT_04 of inst : label is "720D82C8680416B0F0CBF9212F587AF57AA6298E71D9F7A676766674D9C452B0";
    attribute INIT_05 of inst : label is "4930ADABA68CCC97370B24EA15AEE87D0FA16645E743881C424820E17240CEFD";
    attribute INIT_06 of inst : label is "DA54C00AAAA8A02A00080A0AA0A80AAAAAAAA6B65AB20972DDFEDBEB1C192845";
    attribute INIT_07 of inst : label is "31C8F95DA952E90CC54086904CA367A8306EA959B9EA4AF1A8315BC212E344B2";
    attribute INIT_08 of inst : label is "D529B8DE9C8E3CDB7702EE29F241AE80A816D27FADB8E2A4324E6849A229E522";
    attribute INIT_09 of inst : label is "21B06779E71B92823142A552A95480148AB4B4714C2A501250CEA0C360F208A1";
    attribute INIT_0A of inst : label is "4C4E41268508107C7C3F599CBE5985700F2E0B98609F13A058892609C6CC6B8B";
    attribute INIT_0B of inst : label is "304766D8C7080B71999D82154AA2224246E0FB87D89059257E94F8206501624E";
    attribute INIT_0C of inst : label is "0BA04D837007C75C7145145030DC749C74A3E3BF1C03FEDE03F0C5DBF3F3F171";
    attribute INIT_0D of inst : label is "44E82FFD6198BAA282410A34830278D29B6917D719616FCAE058324EB346720F";
    attribute INIT_0E of inst : label is "8F951F7F55AB524F5FE3BFC012218586B8070012A1078B1C1201C74CC605BE7F";
    attribute INIT_0F of inst : label is "AEC002A000B400A8002D8ED6CD6DE9174BE7DF7EF92851551229F8F98F3702F6";
    attribute INIT_10 of inst : label is "C461ED7151701109D97DBD6A959B6FB7AE0CA0F36988C8008404672312D10500";
    attribute INIT_11 of inst : label is "7030079243C818B5BC15022E01D9C94E646589276A63A0ACD26F8D1AB0158C9D";
    attribute INIT_12 of inst : label is "605F8B159687F8441DB9E67CE44DB73619E4550054C4210C434B7B4AD68A6211";
    attribute INIT_13 of inst : label is "DA001907085A3A4A99445A606D367EBCBF8E0B064E79E0CDCEC0F4D99A10B978";
    attribute INIT_14 of inst : label is "0048B5993DDB2467BF61BBBBAEC188ABB24692D4DB5B22288DCD9BB466672328";
    attribute INIT_15 of inst : label is "F3819CC5E7036E9C8CDDA52391FE9CFA71953F4D9AD10153FFF98BD409000120";
    attribute INIT_16 of inst : label is "4C338D83743F15759E3C7392E732C70218E41E62E5CE061C32E61975C357373A";
    attribute INIT_17 of inst : label is "A39206187F8AB693B6A96D5AEB299C61861E3F5DDB58E7593718B9C0CF32E703";
    attribute INIT_18 of inst : label is "2B60769C76E1B7B28B5E28B6CD3745A20A8C795B9A3A8965D96DB61DE5C6D582";
    attribute INIT_19 of inst : label is "844549AEBC68A82340FAE14E0F9DF7294274AC712DCC388CC63108662A7D83D7";
    attribute INIT_1A of inst : label is "20000080FFFCBCDF0000000000A10C4322930642308C623922274E142DE19224";
    attribute INIT_1B of inst : label is "42000000FEFFBD1780000000100A848D00100000BE7FBF7700000000090A003B";
    attribute INIT_1C of inst : label is "EF257386DA72EDEE1E7CCF669A098E624B19A93A68749CDA2C3074D75B753334";
    attribute INIT_1D of inst : label is "55555524A6FE7E7E2FEEDFB399DE608058B13003E162D64FAF7AF521D89A0654";
    attribute INIT_1E of inst : label is "F38E1222E49651DECB9B8D9B6FAD58B6FB938D1FF0CCA0B791747A6B33257654";
    attribute INIT_1F of inst : label is "509DED52E0EF54B60000000804000000F544A220CE99C9860000000600010000";
    attribute INIT_20 of inst : label is "651A8D489203098301DCC5603865300CA01A5D4004144145416D0CB5D633270C";
    attribute INIT_21 of inst : label is "9B69CE183C0394701B20AF759A6D06C7AD866E20000415FBF9F59BB9B9E1EFAD";
    attribute INIT_22 of inst : label is "5F0017FFFE0D99321293AD4D07F29B52F9F7DFBE4ADE89FFD84A2EBB103333CA";
    attribute INIT_23 of inst : label is "6AB2A8053C4D7F7F107855AAD5D7D009E91F557D5C12833EAABEFA1E8F2E2FC1";
    attribute INIT_24 of inst : label is "BBC0754C2B0505E0A0522D948C6003061800003433DAFFA805700FE0E0001AEA";
    attribute INIT_25 of inst : label is "64080102EA5FBFF40000000004800420B2A40020FCFE577E000000083500AAC2";
    attribute INIT_26 of inst : label is "1A8840403BDF4F5E0000000100000400A8410000B9E7E36F0000000081000000";
    attribute INIT_27 of inst : label is "AF5E76CC3CCF2659B7364EBD7EF5FBF43E74E6728205DEDA7DE2031B608A4082";
    attribute INIT_28 of inst : label is "58381D6ADDE380E2E0CB414500360B2094F28E08A0FAF8A174C551CCC8E4FF92";
    attribute INIT_29 of inst : label is "AA6C9B8C90DE437C02A20005544C709FF883220FF3971E593A0F0CB15489D72D";
    attribute INIT_2A of inst : label is "FB4798CC46553AFD17F499322098EAAA688A696E69D8F41DF1C46093B999E496";
    attribute INIT_2B of inst : label is "7AF0BB390988E8DEFE4C01044445F214C19C1E3B0F1CF2177B1E16EAF65A25AA";
    attribute INIT_2C of inst : label is "08B433CBBFF04259E73E33832DAB47C3D0CBC44A55CBD28C78E49B61D5AD57BF";
    attribute INIT_2D of inst : label is "E6A3E32998D91966499BBD2B1B03B7C81DBE501D42A837CC08DC1D99ECE03DD9";
    attribute INIT_2E of inst : label is "EF5A71910CEAFE59D6A275F4141B5FA4252524313453EBBCC73ED31CFB439C39";
    attribute INIT_2F of inst : label is "509CA550E0EF54A60000000804000000F546A2208E91C90612B978CAB0ADC015";
    attribute INIT_30 of inst : label is "49C2D5ABF1488027E238E298E6F8C36DF13C9E7DF79E7DDD1807162967902092";
    attribute INIT_31 of inst : label is "80040002000000090015445001144155401C10A67EB282B963C6C5C522040092";
    attribute INIT_32 of inst : label is "0000004000000000FFFFFFFF9002284B942014040000000077FFFFF7E4005A08";
    attribute INIT_33 of inst : label is "D000800000000000FFFFFFFF75080C477040802100000000FFFFFFFF08B40802";
    attribute INIT_34 of inst : label is "CBD28A58DFFBD7AF00000000400208104EB4502977ADF7EF0000000000000C00";
    attribute INIT_35 of inst : label is "64080102EB5FFFF40000000004800400B2A40020FCFEDFFF0000000002100002";
    attribute INIT_36 of inst : label is "188840407BDF4FDE0000000100000480A8410000B9E7F36F0000000081000000";
    attribute INIT_37 of inst : label is "C24348B4BAF5FAFD000000020000800110B80088FED9FE950000002000002000";
    attribute INIT_38 of inst : label is "10000000DC9F5D7D000000009204000200080020D4BB7E680000004000A06024";
    attribute INIT_39 of inst : label is "0000010035FBE0DB000000004702009604114110F94CC67600000000202A1229";
    attribute INIT_3A of inst : label is "20000000FFFCB4DF0000000000A90C432D000A41F0FFB1E61000001011246000";
    attribute INIT_3B of inst : label is "D0000000FAFF3D1680080000120A888800000000AC33BF77000008000802003B";
    attribute INIT_3C of inst : label is "E120A1E6F77D07702000020000000404C4EEB5A8F131B5A20800000A00000048";
    attribute INIT_3D of inst : label is "F47E1F9CB816211600008004020001008A819DEAF5D9941E0000000400000020";
    attribute INIT_3E of inst : label is "D38E1220C4964BEA1041000000000800DA185E17FC8918698004100000100010";
    attribute INIT_3F of inst : label is "509DE552E0EF54B60000000804000000F546A2208E91C9060000080600110800";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "54A69249042DC4C0431084B0110203C182C40992592C401150FCFE70C0FFFF0C";
    attribute INIT_01 of inst : label is "992412DB44E22A8A1193348B4400EC8104078870F61EFF0DCBEE42A1458C28C8";
    attribute INIT_02 of inst : label is "B2466A3BB912017A16544DF3AEEA4A00100002921CC184AA11520007A550AFB4";
    attribute INIT_03 of inst : label is "A9C7AD84D958B32B105740C0109210118728E4888203097E03A02BDD6ABE29C7";
    attribute INIT_04 of inst : label is "560000002000D7426281C004244854A15225A1B7B7DE7B7083B8D3F80EA46CBC";
    attribute INIT_05 of inst : label is "481643110EC8DD83988163705B59ECBD9792EC0A6701C60F24282052F1406F38";
    attribute INIT_06 of inst : label is "DAADF0A00000AA80000000AA0A000AAAAAAAB236BDF933E245D2CBAB1019A845";
    attribute INIT_07 of inst : label is "FBCC4001B882C52FEE288742AEE52919F73739B45EF74794842108671A660DB4";
    attribute INIT_08 of inst : label is "264CD8586A54DA596DD340400124140C8DD19C39C4EFD560974C4CE0575C2B31";
    attribute INIT_09 of inst : label is "21203085C57304833DCAAD56AB55402DD03C4556D453960201EDE2DBD4960EE7";
    attribute INIT_0A of inst : label is "5EDC41040116024D60B41E1C309E64620F8DC3186480022C2C89B70D7CCE4188";
    attribute INIT_0B of inst : label is "704664DCE609AF39D18822311888A8025194503E8098203D0CA56C0C4500825C";
    attribute INIT_0C of inst : label is "09824D035003C71C71D55D5430D450B450AD6D3D143EDADA23A1E15233333161";
    attribute INIT_0D of inst : label is "4FAB0BFD691E2AEB81B6C4B3982E75C04950E1E498ECA0E06930B2CC4026C23B";
    attribute INIT_0E of inst : label is "AC657D7D61C2166FBBB7F6F8731D41282C25BB205882C10B000D6B96CC5FAC7D";
    attribute INIT_0F of inst : label is "59E17D5406BC5F5501AF5C408409C96AC1BB269936540E41541300E91E51A290";
    attribute INIT_10 of inst : label is "916D14143423DFB69BC94171C4C961202D067A72CDEB0B01879CDF2F167E0892";
    attribute INIT_11 of inst : label is "AEF4A2E291718AA4B81EF7AD55C8DB0DAB759BD2C8731C314806B43620DB0E99";
    attribute INIT_12 of inst : label is "441D7509E539991D0A52C791131DB6665A76676EE9FE73D9678220A42B7F1FD4";
    attribute INIT_13 of inst : label is "058EC8CA8D7F9AB47AFC2B61E95C5738326550E614AAF7FDCA40444ED210AE71";
    attribute INIT_14 of inst : label is "334A79944AB60FC32F1FDD55757D9B5305F35D5B9297BFD17959D5E62C31764B";
    attribute INIT_15 of inst : label is "DBB5CFC5876B6ADBFBF1D67D52750D9C348C676BD37170303BB5100C3961FEE2";
    attribute INIT_16 of inst : label is "6D1147F183860B00CA142DDCE29CF76BCA46DB5AED8ED449E2E5F371A9C093F4";
    attribute INIT_17 of inst : label is "741CBE2022E03326334C2E6043A88A38A38A46D8195E72F7B2D6B1DAE4ACD76B";
    attribute INIT_18 of inst : label is "451E23CF28DC92B31BAFAFBC86A63E160186229088B589688C8D3319C0A241BE";
    attribute INIT_19 of inst : label is "61D4C08048C5592202C4884944447B1086E9FD1696F52F2AAE978F6C9069C161";
    attribute INIT_1A of inst : label is "12002001E40000001810C9008C00410CFC2A351FE85446108CF2140CAB04B912";
    attribute INIT_1B of inst : label is "1280030210E200004206D44A0004449A82220613202800400610210020411401";
    attribute INIT_1C of inst : label is "A42C71B0CE6059474C358625964CA42ACB3BB972CA3DCC0A1C746A9F37AC73B6";
    attribute INIT_1D of inst : label is "555555F664C666662D4A9D31D19C6220749402511DB886612A54A92390B6624C";
    attribute INIT_1E of inst : label is "63049204901041E19173393E11968B6CD1BB370DEC4B66BDB2AC725AF6352350";
    attribute INIT_1F of inst : label is "9500862C9841022041006581024005B98000002619610804008824084088310D";
    attribute INIT_20 of inst : label is "693088409786940100A2542A1C6534AE84611D0AD604505404592EB1D633A5CF";
    attribute INIT_21 of inst : label is "AAEAF444EB397023C9289FADE9C94CB425A3413FFAA9C398D93BD04A4FD6E95E";
    attribute INIT_22 of inst : label is "0667E6DB6D3DF0E60AAA0049A27083706EC9A64D9E798C965B20A2E7194899A8";
    attribute INIT_23 of inst : label is "806931B24510840107058201201006341460000006696C8011400C6820C0F231";
    attribute INIT_24 of inst : label is "603ACA65D0B07A160C190C044A4AAA4DF3F7DFE18EA000515802F0010A66E501";
    attribute INIT_25 of inst : label is "E0600500E400A00000000000000001080004400083A02A090204000010EB1C1D";
    attribute INIT_26 of inst : label is "E1048003006624808000000002000668401400099200840A6820000340D52008";
    attribute INIT_27 of inst : label is "60A6953D7C610A6913AA552A50A152A604F674E292019CCB882E0363E0CE09A4";
    attribute INIT_28 of inst : label is "90B31264C10B32C0DCCB0E6D879208213664CC1DFD0EE661A4EC36DCFCDC13E0";
    attribute INIT_29 of inst : label is "CE2901C0001C007120AC85555C04B2890001638322A70AF3161745E44C992448";
    attribute INIT_2A of inst : label is "89979DADA254556692744BBB601A002CB9C74F78B79D670BB95EE0DB3D1DC896";
    attribute INIT_2B of inst : label is "50D4E2571321C84B1256239F8FDE132C909353796CDD735339075160669B2594";
    attribute INIT_2C of inst : label is "48B041599DD2A60DE63E33822801966B106368E4A08355C610D2400024489428";
    attribute INIT_2D of inst : label is "5365E16B18CACB76A74882B14D63C2531612B02289FB11ED42928B91C251106B";
    attribute INIT_2E of inst : label is "739E50ECBC54462D00032594041A1520606064616C800193D7FFFF7FFF639E6B";
    attribute INIT_2F of inst : label is "9100C62C9801023401006081024005A98000082611E10804B075641FE8509830";
    attribute INIT_30 of inst : label is "DCBB652C32DCA900C018618400687B6DB1B89E7DF79E7DCD0E07870A2D302490";
    attribute INIT_31 of inst : label is "0000672200000010C040050000510155720828367D4260A16C04F5CB72C09274";
    attribute INIT_32 of inst : label is "2044288800000080D9C62E7721400003010A100000020000E3FBDE7B20056482";
    attribute INIT_33 of inst : label is "80244040204000020327E8930400501B2101001B100000009194B0AF00089680";
    attribute INIT_34 of inst : label is "780004286004400B00008000014A100000086000CB180000000440401E020405";
    attribute INIT_35 of inst : label is "E0600500E500A000000000000000010800044000C3A02A090204000000020889";
    attribute INIT_36 of inst : label is "E1048002006624808000000002010648601400099200840A6820000340D5A008";
    attribute INIT_37 of inst : label is "8045181D981405000000000400000301548110C0104449380001020040049404";
    attribute INIT_38 of inst : label is "50002080A00004000900040040701025E2008488180000000048000408882005";
    attribute INIT_39 of inst : label is "180844320004C00A600100203021000044A2000A80004040C00A480101004002";
    attribute INIT_3A of inst : label is "12000011E0000004081089008C004108E2540010000040088200000680420084";
    attribute INIT_3B of inst : label is "32800302104220004004746A0004400282000613200800400600210000411401";
    attribute INIT_3C of inst : label is "A000400208040300028C02980004058800080000610020C08969201001088A42";
    attribute INIT_3D of inst : label is "E001E480E220000284A0080421105B102410000214020403840003020340024F";
    attribute INIT_3E of inst : label is "6204900480100000C28008C202305D8C4800002020000008500A00840004400F";
    attribute INIT_3F of inst : label is "9100C60C9801022401006481024005A98000002619618804048000084288310D";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "40A92C92441CCCC802028038BB22D798D2D2C38400012B2555E4E174C2E0FF13";
    attribute INIT_01 of inst : label is "624C20D244ABB8E81D6CC98B2E01C8C1F16B042CA594099E988EF49AC548B8E0";
    attribute INIT_02 of inst : label is "AC02A950A93529B56486AA8B5041505E021A000B5BC57448A010082D8582CE4B";
    attribute INIT_03 of inst : label is "6116714A3472B309E150000020A5262A4781254468607D3C20F042D09958D869";
    attribute INIT_04 of inst : label is "0C0482081DF40082141039B3800094284141372373C08236E66FA6382873F8A0";
    attribute INIT_05 of inst : label is "3504B03C2B2B97A1AAA9E2314420AA8450AABC2E099AC2D655A54A1A852A2B94";
    attribute INIT_06 of inst : label is "0DBCC8AAAAAA000000000000A00A0AAAAAA0001D2C98AFC1E3B1DBE320D54288";
    attribute INIT_07 of inst : label is "052E0350208814804C27D42B5B001820450220A0C634682706BA08188E142490";
    attribute INIT_08 of inst : label is "02011124B8B2872484F8B824D5CAC4050711786844068404051342A028200802";
    attribute INIT_09 of inst : label is "00805541A0C80441B5000402010076916A98810D18508F21001586B4200D0887";
    attribute INIT_0A of inst : label is "A12144BDC2403A900E07A01E058064060F81E07C1CD022264102190431296D00";
    attribute INIT_0B of inst : label is "0815C922802011AD6F680C964B20C88B5837003668AEC6B143D4769EA00912A1";
    attribute INIT_0C of inst : label is "09824D0302DA1861869A69A6820986A186BF7F382982DAD07001A850FFFFFD01";
    attribute INIT_0D of inst : label is "20044060011E010411F746B79A2E75D0804871F4986862E2E938B2EC6A3EE23B";
    attribute INIT_0E of inst : label is "F605430D0810110F9B07F4693DD1218E811800004080010800000304C45F8000";
    attribute INIT_0F of inst : label is "20D1D55406B8755501AE74DEBDE9E98A69066CB365ACD4451E430401F1C07101";
    attribute INIT_10 of inst : label is "71C9130F4726E1411A4040105540000003101B0BB16202010255DEFB220E6DB6";
    attribute INIT_11 of inst : label is "8CF98A0C85070219B02201AFDD85973808C58952923515D2D602726500A020C1";
    attribute INIT_12 of inst : label is "E2E1019E78011A90A64E94911112485EF2DDD6A7E50647F7DD5029A429570BBA";
    attribute INIT_13 of inst : label is "022F50F9FCDA0EC8361A5A89C76BB3D9C301AAE00A4B3078280114474D7D27B5";
    attribute INIT_14 of inst : label is "0AB494840A61C1126880343CF040A00CC250B08736061088931369C9098C5DF1";
    attribute INIT_15 of inst : label is "EB2EDBBDF65DB69ECE85DEB4C300598165092D0C4255513938535010A6D82120";
    attribute INIT_16 of inst : label is "0D3B6C2303070F604C386C30E630D65D9AD41EF2CDACBA0F82CEC961E3D096E8";
    attribute INIT_17 of inst : label is "E01F018057CC3682370D6D78C391DB6DF718461C1B1AD685371DB5976E78D65D";
    attribute INIT_18 of inst : label is "FE60665B6AE8BA362B3382B3741244000213000500080066180C37279626D181";
    attribute INIT_19 of inst : label is "4B050C981009A14EE80046C3311DC288088AF9451201A618B48463CAE879DB20";
    attribute INIT_1A of inst : label is "820800001080010A8000122800400080130A007998191405B8709B4080602919";
    attribute INIT_1B of inst : label is "021000201800E838000000800002041010008000800008980410410820000008";
    attribute INIT_1C of inst : label is "8D046C60D88B12B41811430049DBA168FB53252024749A1E9D2484100E8C23A4";
    attribute INIT_1D of inst : label is "555555C403DFFFFFA3428D0D6F79402E8A00A058022A86400810200020804669";
    attribute INIT_1E of inst : label is "E20CAEC02004061E2C40E655B134A608510CC500082102D120894CBCA4BE0BE0";
    attribute INIT_1F of inst : label is "B124201D000330206432A005D002018270810405D08200002419901600005121";
    attribute INIT_20 of inst : label is "6D029149B5907600000204080E54A7C8B5AD952B5AD10045054148A9552A4A51";
    attribute INIT_21 of inst : label is "9C69AC26124A742ADB60848DD909483124A6D3110C411DBEDC31B4D85884E10C";
    attribute INIT_22 of inst : label is "CA6BA6DB6CB5D7E77ACE113586C2489A419B2CD96BD89EF6DA4CA68B0E01BB20";
    attribute INIT_23 of inst : label is "BFAEC1FDD5DFFFFE07D57D555FFD78375FD5D555D07FEFEFEEABA06AAABBAA81";
    attribute INIT_24 of inst : label is "7ABAFF05EEBFB957F04024124BCEE46D72DB6DA1FAAAAAAC77F8AAB5BA07AABE";
    attribute INIT_25 of inst : label is "0000000091000000900052008100988444040080C0812000C801884005EBB01D";
    attribute INIT_26 of inst : label is "0000904078040D122210200B59040250000000006110084344002310A00159CE";
    attribute INIT_27 of inst : label is "6480A139131205105245350A1428408320DB5B4011007BC4000802C090A82092";
    attribute INIT_28 of inst : label is "86820204080832021A09040C86800000808052C2880400341185041636369062";
    attribute INIT_29 of inst : label is "A814C434156055822009055000084AD90110CAC9107A40A36026034000012044";
    attribute INIT_2A of inst : label is "304052B90C44C5E7D606022D00731FAE6065BC53B729DE1CE831506CF6D10806";
    attribute INIT_2B of inst : label is "102159620C25100004A72FCE9E9E80902041A0ADD1539FA0EDD3A82B40880180";
    attribute INIT_2C of inst : label is "E038D312662A540294A8A740241840A025A006825420221AA000000C00000408";
    attribute INIT_2D of inst : label is "B6484A465283C204DC000380587C461FEA30C0212223811532866253109D8A03";
    attribute INIT_2E of inst : label is "6B5EAE9B90D3422112C51000094284000000020100508B8141043524105C63D6";
    attribute INIT_2F of inst : label is "B160241D020330200422A005D002018270810401D08200007761C9F1182A6C11";
    attribute INIT_30 of inst : label is "B23E444009138910180000000004306906001629F5926D4086DF22460E814D26";
    attribute INIT_31 of inst : label is "F86E0BA2108C30290055500000041155595430267D15309538253D244E2E1E2C";
    attribute INIT_32 of inst : label is "D960FF6A0000C080B1802068000000007ADD7824121800080028800300000009";
    attribute INIT_33 of inst : label is "5DEFE7B1680424000081005008002010C34368B5308230808F93040100000002";
    attribute INIT_34 of inst : label is "000400000004A0300020C090888D022200000000500061100240EA8C1D082818";
    attribute INIT_35 of inst : label is "0000000091000000920052008100988400040000C0A12000C801884A20034202";
    attribute INIT_36 of inst : label is "00009040F80405123210200959040250000000006110084344002310A00159CE";
    attribute INIT_37 of inst : label is "000200019111000020820049EA1102CD000000000041801116800008241E8048";
    attribute INIT_38 of inst : label is "800000800800218000800002001000020028110B800000800198402200000001";
    attribute INIT_39 of inst : label is "0A9300004E20000000000403A9080200A0040200404082401040004240020212";
    attribute INIT_3A of inst : label is "800800000080010A800002280000008010000040028000001000440200000060";
    attribute INIT_3B of inst : label is "02100020080040BC000004800002041010008000800008980410418820000000";
    attribute INIT_3C of inst : label is "90021808220138440C4F40890000280470081A88002708000000100400801940";
    attribute INIT_3D of inst : label is "C0230011A850020122430086A000202F410800804934B4001111417B40005080";
    attribute INIT_3E of inst : label is "F20CAEC020000700000202200800000966CA104594A091606008400100800000";
    attribute INIT_3F of inst : label is "B120241D020330200432A005D002018270810001D08200000413901601005021";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "80C924925E5EEEE9044310C1D3A467D2CD8A97A512414A68E9031E810100000B";
    attribute INIT_01 of inst : label is "224EB37277443108212449CDCD539B03DA4F00CCAD950B3B2AADC4F2F3CE7A40";
    attribute INIT_02 of inst : label is "CA9C2614480092366DC486639888503E8860102259D924682440082302011449";
    attribute INIT_03 of inst : label is "23142169E5CD71BD0AB8921020A42423479135007948277C44E242C100804261";
    attribute INIT_04 of inst : label is "A4964BE7E3F9E00009670208000480000061392977C2266A2AA22AB1EF27CFC5";
    attribute INIT_05 of inst : label is "22E5B2CCB02A92B0E6B9291240A598831063154C04C05802C6039823081819B2";
    attribute INIT_06 of inst : label is "615D68202A2A800808200A882A2002288880A4DD8D1A2115C5729AEA0872613C";
    attribute INIT_07 of inst : label is "052CA7F36302A02900C59652DA885062044042252104D14400B30C2626840410";
    attribute INIT_08 of inst : label is "2247F6059DB162000EE0AB776A1004018421310A5756A24EA4B95893002B484B";
    attribute INIT_09 of inst : label is "BE594C479242C124A212954AA55281310FB58925190842E081160E9419449108";
    attribute INIT_0A of inst : label is "C2C26DBE7821C8A05629A01C29001155E62A029952B144F54380DD9391296F27";
    attribute INIT_0B of inst : label is "44BCC9329CB2D0A525280A552A92A77BC95728357029446613B676BF107E0280";
    attribute INIT_0C of inst : label is "7C30FF3804CA024024924924F9E824E124E1E1F8483FFFF02903C801FFFFFC41";
    attribute INIT_0D of inst : label is "040807F94B3F020824B2D481BB06F504A4C2282C02067210809C066158B84F0C";
    attribute INIT_0E of inst : label is "C43E69A48010050FFF003C12D2174F41006038716290052C71E00FBE1E2E0020";
    attribute INIT_0F of inst : label is "A5C00000018000000060A668D68C0C135E24A9A54D397BEAB2A0040D8008A518";
    attribute INIT_10 of inst : label is "314B21254542C3033908C1423B25911828298C8A3524ECE1061F7FFF040C0012";
    attribute INIT_11 of inst : label is "8CD9CAC88544324C024AC8684D0813090FFD0D7108F994412313206209CC5122";
    attribute INIT_12 of inst : label is "D929494AAA219441430F95B0003248CED2192453C38D6FAF9288AA8D694C1155";
    attribute INIT_13 of inst : label is "36C033088336AA21968088040789935B53F9EF80B9DC366029649D5726B026B2";
    attribute INIT_14 of inst : label is "8608B5A45A208DBACD1292944A5243204641B64162C2944F2613391B8B184CC6";
    attribute INIT_15 of inst : label is "922A16B52454B012A8A926B464D44111053108922457A26E243B921121020372";
    attribute INIT_16 of inst : label is "8A2A28021215981D4020485694A69455109D12D69568AB020A95054D225184A6";
    attribute INIT_17 of inst : label is "E7E03FBFAA0CA420243842860A4110410412D454525084A22414AD15082A9454";
    attribute INIT_18 of inst : label is "6D2144D4489023243A0342A1FE168D28B6325088602625F65308A4A39724B53F";
    attribute INIT_19 of inst : label is "BDD718DC66BA231F1A840ED532B75A69908EB965206976BB84A472484D51026A";
    attribute INIT_1A of inst : label is "85108000C0023420180020450000000047068A444021860265606091503526E7";
    attribute INIT_1B of inst : label is "222020886300E05100300128001080082001820880F650800008040802000000";
    attribute INIT_1C of inst : label is "0840452A90CB93BC93E12D5B24D28500AAD2830D924C115654E50820C60E0400";
    attribute INIT_1D of inst : label is "1111110B097FFFFF8800000525394FC14000009215E53F300000000230A084FB";
    attribute INIT_1E of inst : label is "A50646287118261E2E4E6350B955B28B9D265C4208800C01088BC4E0A4B08B08";
    attribute INIT_1F of inst : label is "48D2180FF8645C206B0818084000043068452430C14C14581810C60120060084";
    attribute INIT_20 of inst : label is "42ED66B92D0D2D86035FBED768CB6C1B4212328631BFABAFFAA71B632C647871";
    attribute INIT_21 of inst : label is "955909AD87D6C3D69242A89B13FBD96A696495C45113690486BD255312AC95E9";
    attribute INIT_22 of inst : label is "1304736DB60C3A32A613BF0A70CE34D7892A69535CD1AD34D470E592E88A807F";
    attribute INIT_23 of inst : label is "1004284AAAA20001A0AAAAAAAAAAAD02000080008404100100010A1555555568";
    attribute INIT_24 of inst : label is "854500C8254A84A95ACEE3F1E465030619249278555555562AAC555855C00010";
    attribute INIT_25 of inst : label is "0000000000001068280A860F0800479A00000010000400000084800830000AC2";
    attribute INIT_26 of inst : label is "0000100000104A080000A41A40422135001040012520000210009003611008DC";
    attribute INIT_27 of inst : label is "D884E209D63A581252E8000000000002E34949493C903955DD4892410910EDA6";
    attribute INIT_28 of inst : label is "0EA5C200008AB0A2857C9ABE4DD92F9F3BDD293FF5D416AC099A84929295944C";
    attribute INIT_29 of inst : label is "30C20800A202880842100505012991BB86224EBB092A4C85A4DE4988713C2040";
    attribute INIT_2A of inst : label is "441452A914854555A44952488B52002F42249A90B16ACD46E49149265257B25F";
    attribute INIT_2B of inst : label is "00428DA71243820118C691AD2D2D0531490568A7B0770F69A797601BCB2597C0";
    attribute INIT_2C of inst : label is "223108188CC2C48294B8EF2DB2FC1502820AC1110802C021028B259220000000";
    attribute INIT_2D of inst : label is "00580C6456B32314D840A360406300191000C48B1463221431AAE6551E1922C3";
    attribute INIT_2E of inst : label is "4A5241116A1B07360F0A0143E010000848484841417ABFB1536D954DB6531821";
    attribute INIT_2F of inst : label is "40D21808E8645C016B281808400004306C442430C10C18581B6791CCC0000B81";
    attribute INIT_30 of inst : label is "972E3E200311C248004104210800B0FB0052D6AFFDB2EF40165F02444A44C924";
    attribute INIT_31 of inst : label is "F0B45ECB00AA0400804550004105415550721366EBBD57D600293E0C47000465";
    attribute INIT_32 of inst : label is "FD3EFAD53D8400C04040400680000204BB95EC10B04740028040008A00000000";
    attribute INIT_33 of inst : label is "FCFF811C44881C0A30400A16000010007F697740C20024001609500F00210000";
    attribute INIT_34 of inst : label is "01006000D106E4520000014220072445080000808001E0414010200601906201";
    attribute INIT_35 of inst : label is "0000000000001060080A860F0800479200000010000400000084900821445702";
    attribute INIT_36 of inst : label is "0000100040104A080000A41A40422135001041012420000202009003611088D8";
    attribute INIT_37 of inst : label is "00000010400024014048002C38C0880A000000005050200010001806800C809D";
    attribute INIT_38 of inst : label is "2A60016004000000000885480000800260520821830002020000100000000900";
    attribute INIT_39 of inst : label is "AA0000103100A0490280100208800004250000004202B0004003800680800002";
    attribute INIT_3A of inst : label is "811080004002A0201C0020450000000040000443914800900044108040000000";
    attribute INIT_3B of inst : label is "00204080C000E05100300028001080082011820A80F450800008040800000000";
    attribute INIT_3C of inst : label is "5B822D2669258050100100829011200C243800284825043422808D0320100005";
    attribute INIT_3D of inst : label is "031404043010010900C0010C2100000300380C004D86682704800880042002E4";
    attribute INIT_3E of inst : label is "84064628711020010486000028400001C01024206110400000C0000C0CA00401";
    attribute INIT_3F of inst : label is "40D21808E8645C016B281808400004306C442430C10C10581810C60120060084";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "66B24924A66DC5D42B08C23CBD125989FFFA49365B6C312FFFFDFF51E7F0FF3C";
    attribute INIT_01 of inst : label is "449614BA88CB92F35C4892D33408CE0151A2006A2D450B8DD99E52AC41602BCC";
    attribute INIT_02 of inst : label is "1EE2E573382FAE6D920C433D77770801B79FE6790C8690AA105B6493B198DE92";
    attribute INIT_03 of inst : label is "80049494E44AF1A9155E40C212931218D15DB5FFBD67E42419B920C0C06043CF";
    attribute INIT_04 of inst : label is "322904D31C061FFCF0C0FDF7CC484C993305FF94E3C8CB0802200230CC86D0BA";
    attribute INIT_05 of inst : label is "6C3268AAC4C1C806004B004B2ED4CE19C33940646E13289879FC66CCF7E6C4BC";
    attribute INIT_06 of inst : label is "B758B97F75DF5FF5FF7FF55FD5D55DD77775F7B718F79941DDF6FB6B009DA264";
    attribute INIT_07 of inst : label is "78C46D5C38FC5FE4E210431866633138522F383108460C73821502439090964B";
    attribute INIT_08 of inst : label is "468C984C1C14184927827588000004068C119032432CF12072440E402A016730";
    attribute INIT_09 of inst : label is "6DB0A5D1EB3F808219CFEAE572FD001C9AB8F4B3C402122318E060C2CE720CE4";
    attribute INIT_0A of inst : label is "8C8CDB6187DE36432791A01D110003240664191B339318BC08893309CC842F93";
    attribute INIT_0B of inst : label is "3062248842088F18D8C0372B95CB736C0478B295EF18492113985C40EF81FC4C";
    attribute INIT_0C of inst : label is "3C003F001DA4E18F1CF38E3D36C61C0718BF3F398702DAD3A4CD1932FFFFFF27";
    attribute INIT_0D of inst : label is "80388863280E0C30C082040118043400004020E41808202001100340C0604608";
    attribute INIT_0E of inst : label is "428504131932626F1B37D0D0D201E1EE8D19BB32F9C8D39F32EC630404080B01";
    attribute INIT_0F of inst : label is "D4F0AAAA01042AAA804108030030B024CF16EDB76F685B55F2200178A72028F0";
    attribute INIT_10 of inst : label is "906124B1F08B19BC9091422C80930227C404E070C190D8C00C0C462710F896C9";
    attribute INIT_11 of inst : label is "E60C63E271F18861B8227CAC81DCCD1420CDF1F7587AB321D02585B6E0C71CB9";
    attribute INIT_12 of inst : label is "CC9B3B21069BB37C299BC0300000026459261AE838B0230862664B8C60440C11";
    attribute INIT_13 of inst : label is "130029020000281C006867A4259E0E74371C319254FCE3C4C4C2701D98721CE9";
    attribute INIT_14 of inst : label is "335BBFD0188727E79D4EB2B10ACE39F79304C379C8000310CCC8CBB66673375E";
    attribute INIT_15 of inst : label is "C981084D930201DB110D963131BF0CFC3097674BD363AD77342DCA3CDB219F70";
    attribute INIT_16 of inst : label is "6E1107CB56579D1559122130C210C3020C4EDBDECD8604DB62CDB161917DB210";
    attribute INIT_17 of inst : label is "E7FFBFBFAA9EB696B6582F4A4B308820825A575F5B584209B277B0C084ACE302";
    attribute INIT_18 of inst : label is "3C9C36D862CDBF371B8E30BC5C9E6676038631979F13936F59AEB2694782D5BF";
    attribute INIT_19 of inst : label is "8F8DC988384CF9E0E448F987CBF543350E65DC92A48C3D19DE538DE05A758363";
    attribute INIT_1A of inst : label is "A040000800000000C0C210002DBA0C806AE063C670EF4A3260026EEC31C39201";
    attribute INIT_1B of inst : label is "8008000401042000055084018025088AD0000001000004180C19001180680C28";
    attribute INIT_1C of inst : label is "6D2D79C2CE22C8BF0E2CC776DB5CAC2A5B98DC7B6D25DE1C8972261870A172C9";
    attribute INIT_1D of inst : label is "EEEEEE32E41FFFFFE4C99338D894263EBFB9FEB134228723264C9971839663FE";
    attribute INIT_1E of inst : label is "F0481000704001E18B39BC133B06FDE6BB99A48A264F65670626322632132130";
    attribute INIT_1F of inst : label is "FA020001E0A01801E320A0E4065E4580F8000000801204020152000798849322";
    attribute INIT_20 of inst : label is "65BACD6DB60604830188D0683275354EA1029D40000154055575CEB9D73B878E";
    attribute INIT_21 of inst : label is "D96D8CCCF666D0F39B68A7589BE82C63AD92E76AB2A9F5BAD8C1B9C808A6C60E";
    attribute INIT_22 of inst : label is "641C400000882040840441FD0273C333C5BB6DDBCAD89FB6DF80B6DBB9639162";
    attribute INIT_23 of inst : label is "4551400A2A28AAAA00AA8AAAAAAAA808AAAA2AAA281155545554501555545540";
    attribute INIT_24 of inst : label is "95452A80254284A850783C9E00855008216DB640555555502AA0554055015545";
    attribute INIT_25 of inst : label is "A0800680A0C040200000000030300200F000480082800C200000042042144002";
    attribute INIT_26 of inst : label is "08020010050C340000000200004004810000011210000144100008024030C102";
    attribute INIT_27 of inst : label is "FCFE3B6C9CED02690BB243264C99326626B636208A01940823660B22E0CE16CB";
    attribute INIT_28 of inst : label is "9798A44C99797C5E72D3296994361B6C4632C60A00D659E4346073CCECEC845A";
    attribute INIT_29 of inst : label is "CE3DF7FF5DFD77F7BDEFCFFFFC1475939C0B258B35831E11B2072C209C8A4489";
    attribute INIT_2A of inst : label is "BBF38C1CAA156C589624393A6038005099CF684239C17408B2CE20998D8D6136";
    attribute INIT_2B of inst : label is "4C9D72511D02EC487E3795A000019A1C9C9F3B189D1D313318B7326AE6184D88";
    attribute INIT_2C of inst : label is "20302142626C724C624618CB4C83E2F97DF93EEEF7F13FDEFC749A4064891326";
    attribute INIT_2D of inst : label is "6AF663190D0918EE790BA3692B208AC904567001E33910E0880F9781C0C31359";
    attribute INIT_2E of inst : label is "6B5B1391605ADF7930F5FCBC1F89932C2C2C26272CD44B5789043E2410F08508";
    attribute INIT_2F of inst : label is "CA02000128A01801A330A0E406564500F800000080134482DAE05E4230FFF0D1";
    attribute INIT_30 of inst : label is "4186858121C8A000700000000032EB6D9D091E79F79E7DC65D306489E13012C9";
    attribute INIT_31 of inst : label is "C004000400008810C0FEBBEFFEBAAAAAA6E810344BB190B96114618722D4C110";
    attribute INIT_32 of inst : label is "101C6100201000007E87E70A3A7E05044000A00650000000B4D8DB7F9CC0288D";
    attribute INIT_33 of inst : label is "812000000000C008413F32F7317444002000000100100200B457CDCF10E43008";
    attribute INIT_34 of inst : label is "F010000010CC428000092002018400A0D0100400606028000002200184002001";
    attribute INIT_35 of inst : label is "A0800600A040E0000000000020300200F000480682800C20000004204E88A000";
    attribute INIT_36 of inst : label is "08020010050C360000000200004004810000011290000144100008024030C102";
    attribute INIT_37 of inst : label is "F400801046420830000000001130000818010008B0700209002040001C810400";
    attribute INIT_38 of inst : label is "B0000124200000004800200602092A0420014040000000000829128136840A00";
    attribute INIT_39 of inst : label is "70040022200200000041040F9382000412000400400202200001422C6C898001";
    attribute INIT_3A of inst : label is "8040000800000000808000100930008060400086800000041182C40004410A00";
    attribute INIT_3B of inst : label is "8000000000002000051084018020008AD0000001000004180C19000180280C68";
    attribute INIT_3C of inst : label is "C003001A00B80600A0026802849715001010205C804000000120C08440C2CB02";
    attribute INIT_3D of inst : label is "7020001C400140082030800F8A202A9070002019D010000000000200951A0306";
    attribute INIT_3E of inst : label is "60481100704000104990B90201001C411002802021040103C0086548A4284C0C";
    attribute INIT_3F of inst : label is "CA02000128801801A320A0E4065E4500F8000000801244024152000780841322";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "42A00000163484802A0A82A094024901FFFA01365924102FFFF1FE01E7F0FF6A";
    attribute INIT_01 of inst : label is "00060ABCCCCA5281500000CB14094605D086006228450313C88AC025018031C4";
    attribute INIT_02 of inst : label is "4A404021182FAE2CA05CC1102222080030001650088A01E8011B6DB391089A00";
    attribute INIT_03 of inst : label is "00041090E04871A9000C018030B13131915CB0DEF9E3E028009B208040205145";
    attribute INIT_04 of inst : label is "2000000000000002D25800000C40C081022DBD18A1804C2802200220CD06C203";
    attribute INIT_05 of inst : label is "242248A28000810400060002BED404308610085044022910200002C00002C024";
    attribute INIT_06 of inst : label is "920090808A0000A00A2A000AAAAAA0A0A0A0B21108551940549A69A90015E12C";
    attribute INIT_07 of inst : label is "6004440510004004E648031420C32110422F1011084204600017020140899249";
    attribute INIT_08 of inst : label is "26482048040020492602C0000000060380480202031073002008050000294600";
    attribute INIT_09 of inst : label is "209081912A2A8600188889542255B608102850A2800212012080C186C4400C40";
    attribute INIT_0A of inst : label is "88884920000002402611A01C11000124062409193383009C0180040008000E00";
    attribute INIT_0B of inst : label is "2020001008011D0848402221108A20080460A285601800041380504000000048";
    attribute INIT_0C of inst : label is "3FBE3FBB301441041041051032CC340D34BF3F3B4C02DAD624C1018233333029";
    attribute INIT_0D of inst : label is "4F624BFC288E98208375CEB69BEA3DD2926955D6F96D6AEAEF6FB3ACBA5EA7F7";
    attribute INIT_0E of inst : label is "409004100102826F1B7411D0D20164EE9D1BBB3EB949D2973EECEF9ECFD79B7B";
    attribute INIT_0F of inst : label is "5420AAAA02082AAA80820000000000C0C732C5162B400B00F0200128A31028C0";
    attribute INIT_10 of inst : label is "00412DA0A1CBC8B411897C2480010120040C40C0410008000404C46200A1925B";
    attribute INIT_11 of inst : label is "064CE2E431739044942834A4E4AD85B08444D1E22868A32180210DCAD0020891";
    attribute INIT_12 of inst : label is "45921261048A2128613700A0000000041032E6BBB386B40B2F8C0B0840000411";
    attribute INIT_13 of inst : label is "11C621C0630020148228258422B200702518113010B581040042E0100AD600E3";
    attribute INIT_14 of inst : label is "110B2960100522A490442020008411569184616848605130448052124252111E";
    attribute INIT_15 of inst : label is "5B01084CB602014B130CB4202847181C6056650943E1A04E046E862811209670";
    attribute INIT_16 of inst : label is "241107C95452D0150912233242126602084C494A448C044B264D9324B16D1212";
    attribute INIT_17 of inst : label is "100000002A9692869270260A09208820824A124B4948422092D3918085E64602";
    attribute INIT_18 of inst : label is "19B4228C2244951209182098B9842254010620100091016B48A692410D025480";
    attribute INIT_19 of inst : label is "8E848902200450C00044E1860AE010358504CAAAAD883188956A314052248142";
    attribute INIT_1A of inst : label is "00000000E300400505000010D8BBDEF788E023C230E50E22602066F821C10221";
    attribute INIT_1B of inst : label is "100004002220045002000404BDB74FBF000000003C04908008480102F5DBE7BF";
    attribute INIT_1C of inst : label is "450D29424C4681380A0841524908C4701910F5692521CA0C0823220820806249";
    attribute INIT_1D of inst : label is "05050502C0066666040C102848100000008000B13420130020408111149C63F2";
    attribute INIT_1E of inst : label is "0A0000020000061F0A28951122073542220A8882064FC5270202006220110110";
    attribute INIT_1F of inst : label is "12000000080080002F3DECF7146005270400000000000001CABCC1F784F745BF";
    attribute INIT_20 of inst : label is "30985C249302A003018AD56031451428A1085142109455500035A8B516A22608";
    attribute INIT_21 of inst : label is "4D24C468543480F10928AC108A8024430492562AB2A88C964884958908A24427";
    attribute INIT_22 of inst : label is "80008000011040810860008820010071CCB1458ACA488B924FFF125999430042";
    attribute INIT_23 of inst : label is "4551700A2A28AAAB10AA8AAAAAAAAE08AAAA2AAA2E11555455545C1555545570";
    attribute INIT_24 of inst : label is "95452AE43542C6A85C20108841055E30C0000084555555512AA2554455615545";
    attribute INIT_25 of inst : label is "04000000F800402038180107CD9D9FFF000000004044000000E1A005D2145C42";
    attribute INIT_26 of inst : label is "00000000A000002004209222EFFDF7DF000000000980040C00201101B7ECFFF9";
    attribute INIT_27 of inst : label is "98343B2894AC02600EB2402040810206029212001801100829440A2240C4165B";
    attribute INIT_28 of inst : label is "9098A2448969485A624921249092082052965242AA51116010042284A4AC0400";
    attribute INIT_29 of inst : label is "C4000000000000000000055558103582940A018215021C0180042800180A2648";
    attribute INIT_2A of inst : label is "80020008E01508509244102040101F80B1492102205150808288000A84842C16";
    attribute INIT_2B of inst : label is "409520031C0380205C1595A4040580081C9F10088914911148A5122682C80584";
    attribute INIT_2C of inst : label is "0020000666202040000C0A494480120100090000000900000040000024081020";
    attribute INIT_2D of inst : label is "60920208041110447002A00C0220808904046010C1111082080C9401008B1011";
    attribute INIT_2E of inst : label is "210A138060089751000004800048102028202229388001060104180410708508";
    attribute INIT_2F of inst : label is "12000000080080002F05A4FF147005270400000004000001D8A09E42308018D0";
    attribute INIT_30 of inst : label is "810610A100802DB6533EEB9CE62A8B6D94001E79F79E7DC550850649402012D9";
    attribute INIT_31 of inst : label is "FBDFFF7D93040810000100415015544476E000144A31121D2114050200D4C520";
    attribute INIT_32 of inst : label is "FFFFFFFFD21000802020884000000000FFEBFFFF860410180C00006800000000";
    attribute INIT_33 of inst : label is "FFFFFF7F20C1280902490000000000007FDFEFFF189520104200000000000000";
    attribute INIT_34 of inst : label is "080000000200001080E50CABADFFFDEF00001000500400007098098CFC9FE777";
    attribute INIT_35 of inst : label is "04000000F020400038580147CFDD9FFF00000000C044000080C1A005DF2FFDFF";
    attribute INIT_36 of inst : label is "00000000A000002004009202FFFDF7DF000000000800040C00201101B7ECFFFF";
    attribute INIT_37 of inst : label is "0000000003000080090C1233FE93DBAF000000000180000040140105F8DF7CF7";
    attribute INIT_38 of inst : label is "000000008A004A280000020059751D56000000040000000084010000CAF55D65";
    attribute INIT_39 of inst : label is "0000000050240000000000021075E77E00000000100088100001008051EB87DD";
    attribute INIT_3A of inst : label is "00000000C30000050500001048B1DEF38000022080421040044000024A1D29DF";
    attribute INIT_3B of inst : label is "000004002220045002000404BDB30F9F00000000380410800848010244D3C7B5";
    attribute INIT_3C of inst : label is "00008000100000005CC9490157C5F936C0000000200000003DBDE9C2D60B4A10";
    attribute INIT_3D of inst : label is "18000028000000009221AA9C8114E09F80401000000020204CC2642BC101D506";
    attribute INIT_3E of inst : label is "08000002000000000CA0A6A8BBF8EF778000000020000000190AC4417DFF29F5";
    attribute INIT_3F of inst : label is "12000000080080002F35A4FF147005270400000004000001C8B8413784F745BF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
