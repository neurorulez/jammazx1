-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_8R is
port (
	CLK  : in  std_logic;
	ENA  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_8R is

	signal rom_addr : std_logic_vector(12 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(12 downto 0) <= ADDR;
	end process;

	ROM_8R_0 : RAMB16_S2
	generic map (
		INIT_00 => x"04410136040710140605254405D86840FFFFFFFFFFFFFFFF0000000000000000",
		INIT_01 => x"0DC1A46213C81666000024A5000046A0FED040403B9260808208B5902001482A",
		INIT_02 => x"0114510501D190144605254405D8684020A6DFF0D40B3843E0BC6FFDFFFD6867",
		INIT_03 => x"FCFFFCFF3FCF3FCFFF3FFFFFCFFFFFFF020055080002F7FF04004B9E000BFF92",
		INIT_04 => x"FFFFFFFFF3FCF3FCFD7F4113F3FCFFFF0000555520005555FF3FFF3FCFFFCFFF",
		INIT_05 => x"F3FCF3FCFF3FFF3FF3FCFFFFFF3FFFFFCFFFCFFFFFFFFFFFFFFF0010F5FF5013",
		INIT_06 => x"0FFC0FFC0FF30FF30FFC00000FF300FF0000FFFFABFFFFFFFCFFFFFF3FCFFFFF",
		INIT_07 => x"0000FFFF0000FA800FFC0FFC0FFC0FFC0FFC00000FFC00000000FFFF0000FFFF",
		INIT_08 => x"2200EFBE00009FAAFFFCFFFC0FFC0FFCFFFC00000FFC0000F560FFFF0000FFFF",
		INIT_09 => x"E08000C102030107A4890048C89B04410000AAAA0000AAAA0000AAAA0028AAAA",
		INIT_0A => x"2000100140002404DB084021E828008880000088000080230401000400830043",
		INIT_0B => x"001012000018800092802000D2088000008009C02008100040030500C04000E0",
		INIT_0C => x"5810880200800300052104200421000179F10308E2000000E000000002003000",
		INIT_0D => x"4220400A0008008004800020410200023DF400049FF702046048006002004800",
		INIT_0E => x"90A6440812080A120100020048490000F7CF80004B4F000021400C0068208408",
		INIT_0F => x"24082000202021001420080040800800D9FF00014DFEA1001608040000004048",
		INIT_10 => x"01145105011190144605254405D8684043D30000F4F4008081A220210C238012",
		INIT_11 => x"05112D24018DD0F0444187CD0C04C24C0605054405D868405041511604071014",
		INIT_12 => x"FFFFDB73FFFFCD7F0F7DB3D7FDD0090E440187CD0100C24C054609270494B8B4",
		INIT_13 => x"2AAA2AAA2AAA2AAA0000000000000000FFFFFFFFFFFFFFFFFFFFE67AFFFF2DFF",
		INIT_14 => x"1140154055540001ABD5EABF7EAFF77EB041EAB59E9E502A0000000000000000",
		INIT_15 => x"C484C484848F848FFC84FFFF848FFC8F00C300C30C300C3000C300C30C300C30",
		INIT_16 => x"E5A5E5A555555555E5A5E5A555555555010101010101010101010101010F010F",
		INIT_17 => x"C32BC02AFEEFAAAF00FF00FFFFFFFFFF32FF00FFFFFFFFFF00000000002F001F",
		INIT_18 => x"0300FFFE0000FFFF0000FBFF0003000F00000000000300030000000000000000",
		INIT_19 => x"C000FFFF00038003000000000000000000000000000000000300030000000000",
		INIT_1A => x"0300FFFF0300FFFF0300FFFF00030003FFFFFDFF00030003C000C00000030003",
		INIT_1B => x"B9B82E376BBF74FF0000FBFB0280FFBF0000F38200008201FFFFFFFFFFFFFFFF",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFF0000000000000000EDA1820080890477",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"FFFFFFFFFFFFFFFFFFFFAAFFFFFFFFFFDB69EFFFAE78FFFF00570AFFFFFD800A",
		INIT_21 => x"0000200C555B0BFF000000000000000A02C0F4F8001F10FF0010AF2FA3FFFFFF",
		INIT_22 => x"80AA531B800864BB002B0000D016026000000000000F00BF0000000003FF2AAA",
		INIT_23 => x"8EE90000B4FA00000080A903C00FFFFF82FFFFFFFFFFFFFF585007EF0000FFF0",
		INIT_24 => x"00000A80000000180088C00013AC000000000000000000000055051550005500",
		INIT_25 => x"500700BDF00001007C00A0FD4002FE800002FFFFFF40FFFF000000000B7B0ADD",
		INIT_26 => x"00009FBC000080000002AA802000FE1505C8F2AB2078640AEA0CFFFF8BFDF800",
		INIT_27 => x"665F59BFFFFFFFFF5555FC0055550000FFE0FFFF0001F81EFFFFFFFFFFE0FFFF",
		INIT_28 => x"8200E7D02020282BFFC0A95028007FFADE3A52E7F200F917ADFD6E3F8282FFFF",
		INIT_29 => x"F85F0155FDFFC4FFF502FFD404000000BFBDDFBFA000EFBE5BDDEE2B4D5FFFFF",
		INIT_2A => x"0F81285D80255E00BBEF7F7B6EE7FC59A7554AAFB79FFFFF02207F7B0200FEFE",
		INIT_2B => x"AFFA7FD54556E8AAA8AA8AAAB8AAA2AA3A2A002F2BFFFFFFBF9A000F008FA3C5",
		INIT_2C => x"AA4AFF404BA902BEFF66E00B000BFFFF02207F7B0200FEFE00AAFD5580220000",
		INIT_2D => x"9F172E5C91E1BE9D82D4FFFF0A8BFFFFFDD726665D4B173051FB7F5F7EFF5749",
		INIT_2E => x"8002AAEDE9A00003F800FFFFBF2FF000FFDF4081F7FD2084A116E750A26A19D5",
		INIT_2F => x"7F7FEDD5EF3E6657FFFEFFFF5EEFFFFF7899AEAA0A22B82AFFEAFFFF9A8EFFEA",
		INIT_30 => x"13FFF0BFFFFFFFFF4FFFFFFFFFFFFFFFDFFF68B85D8093CB57E3592D111589FA",
		INIT_31 => x"3FFF0FC0CC3300F00A8FFFF0FCFF7FFF303F3C2FFFFFFFFF143FD703FFFFFFFF",
		INIT_32 => x"00A400FF4866FFBF00FC00FC34FC33AF03F507FC40330C33000000000C330C33",
		INIT_33 => x"0FDAFFFF8FF7BFC0FFFFFFFFF540C0D7FFFFFFFFFF50FC3FFFFFFFFFFFC7FFF3",
		INIT_34 => x"FFF0ABFF000FF03C540B0000FC0C3C0CFF00FFF8FC0003F07FFFCFFFFD80FFC3",
		INIT_35 => x"C000FFF0FFFF0BFF001FAFFFB9EEFE7FAAAA0000FFF50003200050000001ECEC",
		INIT_36 => x"55FF5D7FFF55D75FFFFFFFFFFFFFFFFFFFF5FFFC555530C3870D07FF7FD787DB",
		INIT_37 => x"4846AFAA4848AAAA00000E000AAA002C0700F5550034555FE000BFFF0002FFFF",
		INIT_38 => x"FD03FCC3CC0CCEA4FCC3FCCCC3CEC3CCF3CCFCFF02A0F3CFFFFFFFFFFCFFFFFF",
		INIT_39 => x"D000CECE0002C0010000FFFF03FFFFFAC3FF43FFF3F3F1F02FFF03FDFC30000C",
		INIT_3A => x"FFFFFFFFF8148000FFFFFFFFFF80FFFF09B242FB2612EB8A911EE7EEF8006000",
		INIT_3B => x"0002D1052218C40181657FFFFBF4A3F0FFFCFFFF81FDF3DBFFFFFFFFC3BEC17D",
		INIT_3C => x"125F9FDDB9EF1000FA44FFFF4842C89949296F7B1892FBA36410FEFF8101EFBD",
		INIT_3D => x"FF40EFFB4192CFFF0080EFBA20109FFFFE64FF40A4BD4848FFFBFFFFF7B9FFFF",
		INIT_3E => x"0226880700887FFFB98C0A2092A610900221FF740020BFFF0400FFEF4002BFBF",
		INIT_3F => x"0000000000000000079A00962E6D62408020FFF008404E6E001641C47D1B0077"
	)
	port map (
		DO   => DATA(1 downto 0),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8R_1 : RAMB16_S2
	generic map (
		INIT_00 => x"00410044444654470019146C31521411FFFFFFFFFFFFFFFF0000000000000000",
		INIT_01 => x"08029BB90261EDB70000F1A700005EA50D5C040817D1921A00003EBA820936D9",
		INIT_02 => x"44040430415151107019146C3152141104B787FAFF81FC46DF7F0FFA9FE06EFF",
		INIT_03 => x"FCFFFCFF3FCF3FCFFF3FAAAACFFFAAAA8058AABF1252FFFF00017FFF00AD484C",
		INIT_04 => x"FFFFFFFFF3FCF3FCFC0FA801F3FCEAAA2060AAAA2250AAAAFF3FFF3FCFFFCFFF",
		INIT_05 => x"F3FCF3FCFF3FFF3FF3FCAAAAFF3F8000CFFFCFFFFFFFFFFFFFFFCAA3F0FF822A",
		INIT_06 => x"0FFC0FFC0FF30FF30FFC77770FF375AA0ABFFFFFFFFFFFFFFCFFAAAA3FCFAAAA",
		INIT_07 => x"A400FFFF0000FFFF0FFC0FFC0FFC0FFC0FFC77770FFC77772000FFFF0000FFFF",
		INIT_08 => x"585DFFFF0A6AFFD5FFFCFFFC0FFC0FFCFFFC77770FFC7777FFAFFFFFAAA8FFFF",
		INIT_09 => x"35038170107700834020408030038011588855559A0255556A1055554850555F",
		INIT_0A => x"6710220947058E22A008000823A00180001408200046814B0600042110051023",
		INIT_0B => x"5171260A14461A19400400802010010280080050000001000100104860048030",
		INIT_0C => x"0412200014119800110A010010418100241C0114140022480440009000020604",
		INIT_0D => x"2414804291100405102040001000000090D2000824C30000200008018000A008",
		INIT_0E => x"118090C04911020880440080210020007867000010942040001001C005A00240",
		INIT_0F => x"00200002040000214200000108010000D1BE00083C9602008212800108100001",
		INIT_10 => x"44040430415151107109146C2052141125250400194000019100400482400002",
		INIT_11 => x"A80220701B0010181A106186000818901019146C315214115101104040445045",
		INIT_12 => x"ED40FEDB46FFE7FF807960C9440818991A1061860008189BA80668719B788E18",
		INIT_13 => x"30A330A330A330A30000000000000000FFFFFFFFFFFFFFFFFFFFDEDBFFFFEFFF",
		INIT_14 => x"8055055040501454557F502F57AAE9AB6FB70005B51140000000000000000000",
		INIT_15 => x"C848C848484F484FFFC8FFFF484FFFCF00000000000000000000000000000000",
		INIT_16 => x"E5A5E5A555555555E5A5E5A555555555000000000000000000000000000F000F",
		INIT_17 => x"C32BC02AFEFFAAAF00FF00FFFFFFFFFF36FF00FFFFFFFFFF00000000001F003F",
		INIT_18 => x"0300FFC0000000000000003F0003000F00000000000300030000000000000000",
		INIT_19 => x"F800FFFF0003F8033FFF3FFFFFFCFFFC3FFF3FFFFFFCFFFC0300030000000000",
		INIT_1A => x"010000000100000001000000000300030000000000030003C000C00000030003",
		INIT_1B => x"511765C07FFF8E7F9091FFFF0A12FFFF0000542200003BAC0000000000000000",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFF000000000000000077EF2F98D9B26387",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"FFFF7FFFFFFFFFFFEBFFBFFFFFFFFFFFEDDBF7FFEFEFFFFF0006FFFFFD5002FF",
		INIT_21 => x"E400EC10000FBFFF0000000000002BFF1F57D01F0AEFDFFFAA60D6FF12FFFFFF",
		INIT_22 => x"0208AAA8005897DE000F0000F8FE007700000000002F0054800000000FFF2AAA",
		INIT_23 => x"FF5F0020401F00000300FFFFC001FFFF2FFFFFFFFFFFFFFF838003F54A207DD0",
		INIT_24 => x"00B803FE0000800F800BF00049200000000000000000000000085FA00000B8A0",
		INIT_25 => x"000200F4400000000C005410AAFF7FE0002FFFFFD050FFFF0000000007FB0F37",
		INIT_26 => x"BE00FFF400000000AA855F77D080FADA0390DFFF16A7C8FFF9DA573F42FCDD00",
		INIT_27 => x"465B7105FFFFFFFFC000FF0000000000FFFAFFFF0034FE01FFFFFFFFFFFEFFFF",
		INIT_28 => x"2225FFFE888EFFFF13BDFCFA431B201F84FF076FFFCAFBA98894C9EF0485FFFF",
		INIT_29 => x"FE030000FE2202FF52AFFFFEC00ACEA869ABBE6AFE00F8AE77B7EDFF7BFFFFFF",
		INIT_2A => x"00AACF7ED46AAFB8EFA36AEEE6EFB9FB8AA2AABFAAFFFFFF6082FBFF1098FFBF",
		INIT_2B => x"EA56F7AF5680DF7C2A2EAE0A2A2AEA83A92300BF8BFFFFFF40455FE0DBFF012B",
		INIT_2C => x"68262E611A4A8000A14400BF00BFFFFF6082FBFF1098FFBFE8FF3EF8F2FE0A80",
		INIT_2D => x"12D2C650A0028B90F800FFFF28BFFFFF9DBA6062AABF1838FEFFF7F7FB79FEFD",
		INIT_2E => x"AE8023BA1AC0A83CFFE0FFFF0288FF8176F710049DA500100200144D184E8988",
		INIT_2F => x"95F7FB7D5157F5DEFFFFFFFFE659FFFFD1A2CAAAFDEEAAA2FFFFFFFFAA2AFFFC",
		INIT_30 => x"0AFFF0FFFFFFFFFF3FFFFFFFFFFFFFFF3B7FD03B30011AFF0443766B60891D7A",
		INIT_31 => x"B5550FCA5433B0F00FF3FF40FFFFBFFF00073C3FFFFFFFFFFFBF7103FFFFFFFF",
		INIT_32 => x"FFFE00FC2229FFF400FC00FC33FC317FF00F0270D6330C33022002200C330C33",
		INIT_33 => x"FDBCFFFF2770FFC0FFFFFFFFEF004C71FFFFFFFFFA00FE1FFFFFFFFFFFC3FFF3",
		INIT_34 => x"FFFBAAAA0F0FB8BC555500007E2C3E2CFF0BF5D7FC0AABF007FFCFFFFFC0FFE0",
		INIT_35 => x"F000FFFC3FFFAFFFFE41FFFFFFFBFFFFFFF5000054000003FC00000000001010",
		INIT_36 => x"FEAA0C3FAAAAC30F0C3F5D7FC30FD75FFF45FFFE5555B0EBF87E00FFB0EBF8BF",
		INIT_37 => x"993DFFFFBD9BFFFFFFFF0F00FFFF003CC000F0880000088FFE00C0FF002FFFC0",
		INIT_38 => x"3483FCC3CC0CC1D0D443C3F4C3CF8288FF3FFFFFC3F0FB6FFFFFFFFFFCFFFFFF",
		INIT_39 => x"C000C10100070000582802AA2BFFAAAA03FF03FFF1F3F0F0FFFF0140FC30000C",
		INIT_3A => x"FFFFFFFFF782E000FFFFFFFFFFF8FFFF811E6C9762DADFEF9067FFFEFABFE2A0",
		INIT_3B => x"8100FE2816FB0A210601FFFE946803F0FFFFFFFFC03FD555FFFFFFFFC014C000",
		INIT_3C => x"88C9DF505DD54084FE64FFFF691ABFBF8126FBFFFBAEFFFFEB26FFFF1810FEF7",
		INIT_3D => x"5411D7550B9E207D1612BF7F0009506FFBFDFFE8EBB74A12FFFFFFFFFFEDFFFF",
		INIT_3E => x"086E08189B524DD9FFFF9FEE3EFEEC8A98A24400210A017F084467FF1212FFD9",
		INIT_3F => x"000000000000000000771EFFDDD7FEE49000F98E0164C8C202FF28945A219200"
	)
	port map (
		DO   => DATA(3 downto 2),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8R_2 : RAMB16_S2
	generic map (
		INIT_00 => x"00520144524464400058015006141910FFFFFFFFFFFFFFFF0000000000000000",
		INIT_01 => x"4200FFDF0004FFFF0000AC0A000075044740EB372380FBFB0040BB6C0853FEB7",
		INIT_02 => x"001D170500400854405805500614191081F84056D7A0FF503FFF0FFC17FFA5FF",
		INIT_03 => x"FCFFFCFF3FCF3FCFFF3FFFFFCFFFFFFF21010FFFE058FFFF2041FFDB6BFD17E7",
		INIT_04 => x"FFFFFFFFF3FCF3FCF40FAAAAF3FCFFFF46E50000BE380000FF3FFF3FCFFFCFFF",
		INIT_05 => x"F3FCF3FCFF3FFF3FF3FCFFFFFF3FEAAACFFFCFFFFFFFFFFFC01FAAABD007AAAB",
		INIT_06 => x"0FFC0FFC0FF30FF30FFC11110FF310FFFFFFFFFFFFFFFFFFFCFFFFFF3FCFFFFF",
		INIT_07 => x"F000FFFF000CFFFF0FFC0FFC0FFC0FFC0FFC11110FFC1111C000FFFF00ABFFFF",
		INIT_08 => x"6941FFFF2858FFFFFFFCFFFC0FFC0FFCFFFC11110FFC1111FFFFFFFFFE85FFFF",
		INIT_09 => x"1C80859C20034107880020128D0704267FE9FFFF6A58FFFF6BEEFFFF1812FFF0",
		INIT_0A => x"4020401000000060214C0210148602008148574180029517C447D44516651C4D",
		INIT_0B => x"080600000000000204000200018000200400D4FD4000C4450204C6500E00501D",
		INIT_0C => x"00000088001242024080020009120006831020000A0002948A68414C688A51E1",
		INIT_0D => x"840808801448810800000080060100403247000009040002882A112518831494",
		INIT_0E => x"440240004092421000000000020400002908200051B00280A239C510A0A6504D",
		INIT_0F => x"0400020000040080004000080002000043409924410048491A063411B2822719",
		INIT_10 => x"001D17050040005440580D700614392200209020010042480125090408268104",
		INIT_11 => x"73670405C7840000A192CC2267993E14005881500614191014504140500460C0",
		INIT_12 => x"D028FFFF008FFFFFA000C1228E481219A192CC2267993E1C3207340C0D1C9401",
		INIT_13 => x"3BB33BB33BB33BB30000000000000000FFFFFFFFFFFFFFFF7F57BFCF77FF9FFF",
		INIT_14 => x"2552005512A25015FFEDDDAAEFFF83E0DAAD0154ED5D01540000000000000000",
		INIT_15 => x"C484C484848F848FFFFCFFFF848FFFFF00C300C30C300C3000C300C30C300C30",
		INIT_16 => x"E5A5E5A555555555E5A5E5A555555555010101010101010101010101010F010F",
		INIT_17 => x"D57BE02AFEEFAAAF00FF80FFFFFFFFFF10FF00FFFFFFFFFF00000000003F002F",
		INIT_18 => x"0300FFC0000000000000003F0003FFFF00000000000300030000000000000000",
		INIT_19 => x"FF80FFFF0003FF83000000000000000000000000000000000300030000000000",
		INIT_1A => x"FFFFFFFFFFFFFFFFFFFFFFFF00030003FFFFFFFF00030003C000C00000030003",
		INIT_1B => x"72B0441B877FFBFF6149FFFF6858FFFF000049EF0004FFF4FFFFFFFFFFFFFFFF",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFF0000000000000000027705DFFD22F5D4",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"FFFF07FFFFFFFFFFAAFFBFFFFFFFFFFF7FE7FFFFB6F9FFFD002EFFFCE800BFFF",
		INIT_21 => x"0000FC0300BFFFFF0000000200005457A0B763047FFF07FFFFFFFFFF7FFFFFFF",
		INIT_22 => x"80685D01AAEBC098000100001D11000A00000000003F0000100000000FFF2AAA",
		INIT_23 => x"40C05400000000000D03FFFF002FFFFFFFFFFFFFFFFFFFFF47F8000080842000",
		INIT_24 => x"005FAAB7E8006ADFE59FD000BA00000000000000000000000AFC11FDBC000798",
		INIT_25 => x"000F00D00000000003ED0000FF4003F5FAFFFFFFFA80FFFF000000000EFD0FFF",
		INIT_26 => x"FF80FC00000000000160F553201AB9EA0045FA5F557A03DBFDFD5540B0700000",
		INIT_27 => x"9ADB6000FFFF0555E000FF8000000000FFFFFFFF8032FF80FFFFFFFFFFFFFFFF",
		INIT_28 => x"6CC9FFFF8BFFFFEFF901FC860000DDFBF58DE1CA599B6AADE220997FA288FFF9",
		INIT_29 => x"7FEF1000FCA447FFE807BDFFE800E9FF7FFB577DDBBBEF7BDD55BFFFFBFFFFFF",
		INIT_2A => x"FD77D5DB577FD6DEFABFFEFD9AEABF6EA0AAABFFAFFFFFFFADB6FFDE6D99F7DF",
		INIT_2B => x"F4FD5F7BD0A857FBA9CA2ABCAAA2A82A0186CBFFBFFFFFFF80286A116554FA04",
		INIT_2C => x"017F55D554519000FE151BFF0BFFFFFFADB6FFFF6D99FFFFFFFFD5FAFBDF3D00",
		INIT_2D => x"E97E886CFD9D14C0FF83FFFF0BFFFFFFDBBF0000FFFF40EABEA2EF7FDBA9BDEF",
		INIT_2E => x"A4A88111014200A4FFFAFFFF055FFFF0664C00009C65000000295518820031EF",
		INIT_2F => x"754FFFDD7FBD5BDDFFFFFFFFFFB8FFFF88ABFAABA2A9AA0AFFFFFFFFFE22FFFF",
		INIT_30 => x"E7FFC3FFFFFFFFFFBFFFFFFFFFFFFFFFF9B1FAA4697814FB0A65772C3B14CA4D",
		INIT_31 => x"00000FCF0293F0F20FF0FC0BFFFFFFFF00033C3FFFFFFFFFFFFF730BFFFFFFFF",
		INIT_32 => x"008200FC26911CE800FC00FC33F03031FC2F03F000330C3303F003F00C330C33",
		INIT_33 => x"DBFCFFFFBBB0FFC0FFFFFFFE35AA0FF1FFFFFFFF0DBFFF0FFFFFFFFFFFE1FFD1",
		INIT_34 => x"FC0FFFFFFFFFFFFC000000003FFC3FFCFFAFF0C30C0FFFF003FF6FFFFFC0CFF0",
		INIT_35 => x"FE00FFFF0F6FFFFFD8AE55551410555500000000AAFF0003FC00000000000000",
		INIT_36 => x"AAAAAEBFAAAAEBAF0C3F0C3FC30FC30FFF00FFFF0000FFFFFF87003FFFFFFFFF",
		INIT_37 => x"FAFF5555F50B555555550F005400003CC38AF0CC28B00CCFFFE0FF5702FFF56F",
		INIT_38 => x"B8C3FCC3CC0CC20CFCC9C3F3C3CFC3CFFFFFFFFFC3F3FF3FFFFFFFFFFEFFFFFF",
		INIT_39 => x"C000C000000000000EBE02A9BC0F7FFF83FFC3FFF0F0F2F0FFFF0333FC10CC0C",
		INIT_3A => x"FFFFFFFFF07DFFFFFFFFFFFFFFFFFFFF80842B8E25FFBFD59EA5FDF0BFD53370",
		INIT_3B => x"A219B86F829FB97CD288E7FC81F003FAFFFFFFFFE0BCC000FFFFFFFFC228C33C",
		INIT_3C => x"1980D450CAA068A3FED1FFFF0062FFFF3960FFFF15EEFFFFB271FFFFB139FFFF",
		INIT_3D => x"4499FFD01FB78008E410B7F492414045FFFFFF44CD409AD8FFFFFFFFFFFFFFFF",
		INIT_3E => x"897917FBF46A2280077519DE7744FF8861A30000CB960000C81100458C929110",
		INIT_3F => x"000000000000000023BD08441010510896082EFF0008D189081679FB7BFBEEE8"
	)
	port map (
		DO   => DATA(5 downto 4),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

	ROM_8R_3 : RAMB16_S2
	generic map (
		INIT_00 => x"0501301D076120410111201310100014FFFFFFFFFFFFFFFF0000000000000000",
		INIT_01 => x"9A0CDC99A602D9FD000096D9000062EE05E0DDFD01419DDD44009DFD1232DDFD",
		INIT_02 => x"1100444004084711C111741310100014FBF880F35FE8BE283FFE07D301BDBD1F",
		INIT_03 => x"FCFFFCFF3FCF3FCF2A8AFFFFA2AFFFFF4841FFFF34B9FFFF018BFD99BBFB9C1B",
		INIT_04 => x"FFFFFFFFF3FCF3FC102AFFFFA8AAFFFF4121FFFF4249FFFFFF3FFF3FCFFFCFFF",
		INIT_05 => x"F3FCF3FCFF3FFF3FA8AAFFFF2A8AFFFFCFFFCFFFFFFFFFFFA000FFFF0002FFFF",
		INIT_06 => x"0FFC0FFC0FF30FF300A855550028555FFFFFFFFFFFFFFFFFAA2AFFFF8AA2FFFF",
		INIT_07 => x"FFA8FFFF0001FFFF0FFC0FFC0FFC0FFC00A8555500A85555F80AFFFFBFFFFFFF",
		INIT_08 => x"49A9FFFFF859FFFCFFFCFFFC0FFC0FFCD0A8555500A85555FFFFFFFFFFFFFFFF",
		INIT_09 => x"A7A20106209B424301110208030600204948000058590000498E00005958003F",
		INIT_0A => x"002E4512282205060120020062108800408080800140001300920001400B8803",
		INIT_0B => x"82829109924804492004A000811209004200200700400880144C080946510043",
		INIT_0C => x"06060C000882201840024000004012001E6C0200005240021006600000500006",
		INIT_0D => x"2610102020A10008040040000000202040302068407204829E10004010520818",
		INIT_0E => x"8221021022018010000001020820080890108204181EC102042000280500020A",
		INIT_0F => x"80210000102004040000000040002088042C4182609442491080100402122108",
		INIT_10 => x"1100EAEF0408ABFAC111FFFF1010FFFF40408060028042920201000109000188",
		INIT_11 => x"93C300006C580400CB6DF7B6E1DFC1620111FBBF1010BEBE0501FBBF0561FAFB",
		INIT_12 => x"FE6DFFFF67BFFFFFCA4CE2B623C7CF63CB6DF7B6E1DFC96390D2900746210400",
		INIT_13 => x"AAABAAABAAABAAAB0000000000000000FFFFFFFFFFFFFFFFD000FFFF17FFFFFF",
		INIT_14 => x"010A5555AA005555FEF54AA155FF5741FEF555FE55FFBD520000000000000000",
		INIT_15 => x"C848C848484F484FFFFFFFFFC84FFFFF00000000000000000000000000000000",
		INIT_16 => x"E5A5FFA555555555E5A5E5A555555555000000000000000000000000000F000F",
		INIT_17 => x"C02AFE2AAAAFAAAF00FFF8FFFFFFFFFF00FF00FFFFFFFFFF00000000002F001F",
		INIT_18 => x"03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000300030000000000000000",
		INIT_19 => x"FFF8FFFF0003FFFB3FFF3FFFFFFCFFFC3FFF3FFFFFFCFFFC0300030000000000",
		INIT_1A => x"000000000000000000000000000300030000400000030003C000C00000030003",
		INIT_1B => x"06EF531998AFDD6F6B6BFFFF42C9FFFF0000DDCF000F05FC0000000000000000",
		INIT_1C => x"0000000000000000FFFFFFFFFFFFFFFF00000000000000000824120277BD4224",
		INIT_1D => x"0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"FFFF03FFFFFFFFFFABFF3FFFFFFFFFFF8FBDAEEBFF7FEEEF00FDAAAB4200FFFF",
		INIT_21 => x"0008FC2F02FFFFFF000000240000000AFD4F040041FF02FF55D5FFFFBFFFFFFF",
		INIT_22 => x"BDAE202267DF0083000000000024000F00000000003F0000000000000FEA0054",
		INIT_23 => x"00380000000000000C01FFFF2BFFFFFFFFFFFFFFFFFFFFFF0FFF0000FFFF0000",
		INIT_24 => x"0000BBAF4020FEBFD00F4000D400000000000000000000000FD502020000F3E0",
		INIT_25 => x"002F3BCAA800800003FF000050002FF4FFEAFFFFA954FFFF0000000103FF1FBE",
		INIT_26 => x"50000000000000000010FFEA7F20AAAA05028A03AF71C7FFFE78000B8010E000",
		INIT_27 => x"1BAF8000FFFF0000F000FFC000000000FFFFFFFFC031FFE0FFFFFFFFFFFFFFFF",
		INIT_28 => x"6F9AFFFFD540FD5456AA5401800055551D92FF55437A55757E7F6B6FEFBFFFFF",
		INIT_29 => x"07FFFA0AE4FF5955FFA36DDF577AC07F8BDEE757AAFBDB6D17BFBFFFBFFFFFFF",
		INIT_2A => x"0AAABF769401B7ED656D6A6B777EA2E6AABABFFFFFFFFFFF9D9E7F79CB7BC65D",
		INIT_2B => x"D6E977F655FFFDFBAA1A2ADAAAAE6AAA024BFFFFFFFFFFFF55F44A52A8212A5B",
		INIT_2C => x"F8002BF5000040000140BFFFBFFFFFFF9D9EFFFFCB7BFFFF51157FD75FFFBEA0",
		INIT_2D => x"556E5EE90B893BA0FFFFFFFFFFFFFFFF9E360000A15500A8EF7D9EA6F7BFB7EB",
		INIT_2E => x"B2EEE000802A284BFFFFFFFF80B5FFF848B1000032610000E9458445B8270708",
		INIT_2F => x"DF9EFFFDEADFF6F7FFFFFFFFFFA9FFFFA9AAFEBEAAF22A2EFFFFFFFFFEB8FFFF",
		INIT_30 => x"F03FC3FFFFFFFFFFFFFFFFFFFFFFFFFFDDB844A5A79F0000EDC48C891B2F08AA",
		INIT_31 => x"A0000FCF00C1FCCBAFF0F03FFFFFFFFF7D7B3C3FFFFFFFFFFF0733FFFFFFFFFF",
		INIT_32 => x"00FE00FCDBED2CF000FCC3FF33D1C0347C3D03F00C330C3303F003F00C330C33",
		INIT_33 => x"BFFEFFFFFFD5FFC0FFFEFFFFC0FFFFF0FFFFFFFFF07FFFCFFFFFFFFFFFF2FFF3",
		INIT_34 => x"57FFFFF5FFFCFFFC0000AA003FFC3FFCFFFFFAEBAC0FFFF08BFFFFFFFFC2CFFC",
		INIT_35 => x"FF80FFFF01BFFFFF7FEE0000248600AAAABF0000FFFF0003F4007771CCCC1113",
		INIT_36 => x"FFFFFFFFFFFFFFFFFFFFAEBFFFFFEBAFFFA8FFFF2082FFFF7FF800077FFDFFFF",
		INIT_37 => x"DFD400000001000002AA0F00AAAA003CEAAAF064AAAA064F7FFEFFAB2FFFF2BF",
		INIT_38 => x"FCC3FCC3CC0CC38CFCCCF3CFC3CD4147FCFFFFFFE3C3FFFFFFFFFFFFFFFFFFFF",
		INIT_39 => x"CCCC4444C0024DDDBFFFC3FFFFF5E157C3FFC2A8F3F053F003FF0133D000CC0C",
		INIT_3A => x"FFFCFFFF0000FD7FFFFFFFFFFFFFFFFF4608F7BD0917F9001EF4F430F4003330",
		INIT_3B => x"109EEEEBF40BFDFFBE7F2FFF83F000FFFFFFFFFFF0F4C33CFFFFFFFFC33CC3BE",
		INIT_3C => x"E7BF89A1BD14A262FFB7FFFFB889FFFFEDBAFFFF4C7FFFFFEFEDFFFFBCE6FFFF",
		INIT_3D => x"69B93C8237FD29B7BB98052289B92060FFF9FA6D0062F9EFFFFFFFFFFFFFFFFF",
		INIT_3E => x"21FF611DFB76749A20088608400044D2B7AF08189EF6202179B9002289A60080",
		INIT_3F => x"00000000000000006D41820800061820E64B077E4000EFFF084001656FFF3445"
	)
	port map (
		DO   => DATA(7 downto 6),
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => "00",
		EN   => ENA,
		SSR  => '0',
		WE   => '0'
	);

end RTL;
