-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cpurom is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cpurom is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FB4D3B69A6C0C04A8D6098C1151AC1318A8D504DBA0850B2D4050007220A0509";
    attribute INIT_01 of inst : label is "8DFFB8E5CAA734412544B9358F8895B139B27B69E6DA46DE6F4D8FDEDB07E9F3";
    attribute INIT_02 of inst : label is "26335B8E4A862419EF8BFFE022B5A24AD461B8BAF2EEBB7A4F95386CE2A2C51D";
    attribute INIT_03 of inst : label is "8884244A21245515EFAA46691269366226655CD20999EB26E6C6641224D81012";
    attribute INIT_04 of inst : label is "85D09840407DDE6EC635DA6C96AAD446B6EBFFD0A4442FAA9415EA020A024228";
    attribute INIT_05 of inst : label is "9B3F51B2936926D26DA55B6DAAE618A459B3D07ABF4B71F0E101DC0B95B60395";
    attribute INIT_06 of inst : label is "5462A31513B8715495FF7B3F7ACF7A3B2FFCACAFF2B37FAC5159FC668AC99F3C";
    attribute INIT_07 of inst : label is "67B330CE64B33BDE7EF6677BCF90AB5DECF1D385079642487BACE97A21B16104";
    attribute INIT_08 of inst : label is "CCCE40D243AFF8CA6A5B65CC65CE399630B3F161A8D9EF35C008000425FFFFE8";
    attribute INIT_09 of inst : label is "FFCBD11B2E3892811AF4DB083D1D4732EE1B81B0AEAE54B50425542013027D09";
    attribute INIT_0A of inst : label is "203C5447FF7DF1E928C3DC9E10A47C1C2EF9E3918A2B267D7B92C94C95B417B4";
    attribute INIT_0B of inst : label is "104E0C1D258419B2127B404878A8FE3EFBE3FACDC7CDCC506E2DC4B8DC5D8243";
    attribute INIT_0C of inst : label is "7AFBA2560CFFE66DABE54478CF7DF7D8C615323C64444612A5A8199F425D0020";
    attribute INIT_0D of inst : label is "398C4A3DB8C6E358E6A5D94B55555A0DB0CB0D98CD8F024BA20532632D692692";
    attribute INIT_0E of inst : label is "23E0E3021B842A8208B0548ECA912A8208A604FE92692488E79F9F9C67762AE4";
    attribute INIT_0F of inst : label is "3971D49259E6240000014E80850B7552C891CA7DBD51B56F7C49547D5E87FF1F";
    attribute INIT_10 of inst : label is "096A8C64D76552ECFCF54D445734AB21015AD37CFA670DC55BC5FA49FA41FB6E";
    attribute INIT_11 of inst : label is "0002000801100003D13E91F4999D9A82A4A82A4880D00D4E12A844BB94158857";
    attribute INIT_12 of inst : label is "2E4050DC0702449815409B86D2804546ECDC1D080A0DB5484A909A2552242391";
    attribute INIT_13 of inst : label is "936DF74BAF5DCCE556590D8654D14496655540526A34AE6582A62758A8304548";
    attribute INIT_14 of inst : label is "57FC1687F8D7146BF1FC4A8478C7151C580670438E8478C7998A122A52D083DD";
    attribute INIT_15 of inst : label is "87806910357B80F512A10E079B96C0F7EFFF930AFE5CB9457F50A4DB7E387FFD";
    attribute INIT_16 of inst : label is "6722984C2315B82468F718DC5E11556DBF307FE1EAB1BFD29F2F8A487F336596";
    attribute INIT_17 of inst : label is "3B64CED927B7C67228B4292ED906ED914D38016481F4EDDF45F7A154C356A8FF";
    attribute INIT_18 of inst : label is "EBC235D9A8692805E177DCCE7307546D0E4EFF22B951DB20DF7B22D36987F364";
    attribute INIT_19 of inst : label is "011650008ADDB3FE444216AB3094F18B8670C210B92BFB69BF4B84AA44D38756";
    attribute INIT_1A of inst : label is "100E5FAB059D68D7CC8AD281412AB649D612C93A80657A001C6E7F3CE78F3CA0";
    attribute INIT_1B of inst : label is "7AD753861929033552500A997A5F8D5C5D5C521084CF202014A437443291C692";
    attribute INIT_1C of inst : label is "5A06F3C910010912609C8846929EAE79FFDFFB8452528A8ACAC8A2A2A2A26198";
    attribute INIT_1D of inst : label is "66966DB1D1E4198109A130779F981F61D0D098C86B990C93FDC4AFA1327099C5";
    attribute INIT_1E of inst : label is "535C3B2A0A514F3B8FD3C40E7EB7E99C54045D0B0215088A55B3D868529A4964";
    attribute INIT_1F of inst : label is "5E911FCFF53152B0A299131118807A6B9C69068B4CFB62A62D16ABD746CC205A";
    attribute INIT_20 of inst : label is "5F653B2E79609EF2DFE930C0F9660AE20246108F47FFEA791FFD4D5E9E3FFF52";
    attribute INIT_21 of inst : label is "8C16AA2C6AA215E3300236A90A68254060A140CFE5844410CFFFE9F831A24C32";
    attribute INIT_22 of inst : label is "3D19D32360E32601A8C4ACA59124EAD28C738000305510180075900134020026";
    attribute INIT_23 of inst : label is "00000000006060404021010000202121416141202160406AA6DF53438675E19D";
    attribute INIT_24 of inst : label is "080004A00010000AAAAAAAAAAAAAAAA440000000000000000000000000000000";
    attribute INIT_25 of inst : label is "976646046C7A1D6907882622350F3FEC6FD55B7DFFFFE03E0080540C55D40C08";
    attribute INIT_26 of inst : label is "3AA91AD5A748998D0AA9CD014405183B800C94E1171A7175267318C08D08F04A";
    attribute INIT_27 of inst : label is "2EA4B0A0A79AB4E81331A15538D1A740998C0829C68D38998C082DC5B71352A6";
    attribute INIT_28 of inst : label is "D389297525A5453CD9D6E3E97A712C0456F2D829D96E692598F2555B8F1A7125";
    attribute INIT_29 of inst : label is "B689F649936EDA27DB5B71331A1552891B7593318105225E3671652585159E7A";
    attribute INIT_2A of inst : label is "535E8930CC318CEB186B277D3EDDDBFE28BCA19A363F6CC91E5967CF2CB9659F";
    attribute INIT_2B of inst : label is "1111110000000011111111111111117E8398404413EDB6FDACD340C926837095";
    attribute INIT_2C of inst : label is "5F55FC04402000001666667DD50550544150A0082A0A20008A0AAAA88A820911";
    attribute INIT_2D of inst : label is "2222222222222220000000022222222222222222222222311501454150146A91";
    attribute INIT_2E of inst : label is "0055011015011405041104110411500044441044104410462220404222222222";
    attribute INIT_2F of inst : label is "0A280882202880008AA088A0005022288D880202502225401555555050510511";
    attribute INIT_30 of inst : label is "B70AD7FF05550554550554155411677AFDFF8FF8FDFEF9BEFE9EF9AF23200112";
    attribute INIT_31 of inst : label is "F704143A01015151CDD051455054554044446622455514505010000040010541";
    attribute INIT_32 of inst : label is "6AA2582903011105141567313330333311EEFDFCFD6515545155515415500010";
    attribute INIT_33 of inst : label is "D68D02B5017555555055551551DDC98100111015541572275554555511011550";
    attribute INIT_34 of inst : label is "00000000277775DDDDCFFF777731677BFDFFDFF8FFFEF9BFFFDFFDFFFFEFFFFF";
    attribute INIT_35 of inst : label is "00000000000000000000000000000000B1834E09EA4E456D705F7EFDF84A2644";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "5202E6EE66939474AA7653B24034C0D30D30D30D30D3FFFF1D88F26FACE0DFF9";
    attribute INIT_39 of inst : label is "0BEF817D3F0FC0BF7E1C4E0458C0D2ABA02827E0936F6426DEC84A7653B2F9C1";
    attribute INIT_3A of inst : label is "0C6575D1E3E222AF68DEC550921362B3E6AC9C3564F2926949269000B49310B0";
    attribute INIT_3B of inst : label is "9A696A41000A50017E2000C10BC0FCAFF8176B741209FD53B2092906417FAFD0";
    attribute INIT_3C of inst : label is "BE6B5E35AF9AD78F6BE6B5F7DBEFBAD75BA5B1F96597ADD2D8324AB26B2CAAC4";
    attribute INIT_3D of inst : label is "8ACDB0833D65936B1F35AF9ED78D6ABD8F97B5E3DAF9ED78D6BC6B56D9AD78D6";
    attribute INIT_3E of inst : label is "000000000000000000000000000000006DECD3A3EDBE133B25C4B76640406607";
    attribute INIT_3F of inst : label is "0600000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "8CB3068A215C2688460B33CA642C92279AC8A24C88A28400FA0100034C330181";
    attribute INIT_01 of inst : label is "130069113459A75157230642634D1AC64067AFFEE9C85F412DA5C201E54232A3";
    attribute INIT_02 of inst : label is "11090728099D049B4A1DD513ECE8677C32C6155D74B557AA805A468008C9F93B";
    attribute INIT_03 of inst : label is "7556BAAB67BEF3BD46532FACB4704B4D8017B7F4774AA01283DD2CEF6D12DD9F";
    attribute INIT_04 of inst : label is "63451F7D948960016A9A84891C3A467C544500294B0A47A42CFBA64E4E5D556D";
    attribute INIT_05 of inst : label is "49A90D00095C12B800BE00057017247CA2CE3C9726E20DE7A8BC31B795A69D2B";
    attribute INIT_06 of inst : label is "888DCCAA27D745A7FB34C8E4C994C4555911357444D41149EE6E8A4911500450";
    attribute INIT_07 of inst : label is "9864EE119365E413817CBC82711B95A243FA2648E1DCD40DC0AE30DC7EDD6C68";
    attribute INIT_08 of inst : label is "BB9F2F9FE679B799B5F6CB5BCB59EF2DEC6C8B72428054068D9122773E04020F";
    attribute INIT_09 of inst : label is "450664D00147EEA8B8999B6372F137EE6B36F36F1B18FBE6FF4FAB811A503273";
    attribute INIT_0A of inst : label is "3C829980B6C96224B42631393B40C1B279A4DE6D3455401AC44924924A892EFB";
    attribute INIT_0B of inst : label is "6ECF4D61FE4ED5F0A1806F9105732C0D92C42FD560888924DBE44981B7C70D0C";
    attribute INIT_0C of inst : label is "B5CC7EBFC01F4C07258998B756C96C95268702E1A999DA7EF2BC800C9682DC96";
    attribute INIT_0D of inst : label is "6DB4AD458D88EC6D2C632B62BFAFA93E13A80CCB8EECA33C44628C9ABDA5DA54";
    attribute INIT_0E of inst : label is "41685C9E34002ECEEDC3987B58156CCCCD44B9525DA54893004D3236AD96C692";
    attribute INIT_0F of inst : label is "444A6F8CD05A52CADA2B80C69CCEC4DD8CBFE58304C2B76EC08080846A0A800B";
    attribute INIT_10 of inst : label is "F7BB2B5C4968CBA9919498D6DF62C4A4933D9E31CC012DA87FE21EE00AC30612";
    attribute INIT_11 of inst : label is "67A44A7B33F9129B99F5D7AEA99DD8799E47B9ECB312C50DEFA644911A260846";
    attribute INIT_12 of inst : label is "AC0CC4A0B81B9DD26009949CEB338DC52CA4D4672B8A7667E44A7B33F9129BD6";
    attribute INIT_13 of inst : label is "BB6DE00248168346C49681CF32BA4B68197FDCC5ADBDC81804F0EA6B01412365";
    attribute INIT_14 of inst : label is "FFFF379C0E80983C10C2B6117BEF3F94FFEC96DBEA117BEF28811C0D7EBA9A80";
    attribute INIT_15 of inst : label is "34FF204D9103A4A1F1BEDBF81FC7AD891070AA780F3E7CEC07E56EDB7B4D0401";
    attribute INIT_16 of inst : label is "1EE5FCFE7F3DF9862F0072DA3EA31C97280AFADFFC0102012AC54516810076D9";
    attribute INIT_17 of inst : label is "0DBB412A4438601F9D8FBEF65CA34D8AB2022291CC0EEEB06FE0124E015CEA41";
    attribute INIT_18 of inst : label is "B558FAA366C3414EA478249089DC3898B7B00024C01ECB946963152D70300000";
    attribute INIT_19 of inst : label is "68BA85B45487C1F5669921F43D31117CD41754B11D40BEC00BFB1FEFB7E769A8";
    attribute INIT_1A of inst : label is "395F8166FF3B6C0083A28BD39C4FA2E0488E05CE1D9C9DBAB031108510A0870B";
    attribute INIT_1B of inst : label is "80B8E0BAA3BFA46C86829CA9B00238888897EF7FFB9FC4F78F7EBEB7BBFB0CFF";
    attribute INIT_1C of inst : label is "AAA10801A9E7E0400670DE2CFF71F1060020804E9FEF35137151CCCD44454804";
    attribute INIT_1D of inst : label is "2749AA483ABEC04CB6925E18E0128073A9C1DB00E790200100A7F0BA046D034F";
    attribute INIT_1E of inst : label is "8035E4D67D6522092C000BFD98021260E4B979EC99306490EF01BDACE34C9723";
    attribute INIT_1F of inst : label is "346C8582C24CAD67C92D2CE9B346F8066336E6528E53ECF7BBE10032093149AA";
    attribute INIT_20 of inst : label is "CE007005B66D246D8302CCCD621DD67670208A9E216D84B885B0923E050B6C24";
    attribute INIT_21 of inst : label is "C8C0CC680CC60300D00755F89241C00581C4070875B1F6E33207649EFBA48D04";
    attribute INIT_22 of inst : label is "0929951500A01504B42118E6880E4B60880400005866080000439003AE620075";
    attribute INIT_23 of inst : label is "454545454020202021E1E1E1E1E1C0C0416141A1A061200CC9CD0583CA64C299";
    attribute INIT_24 of inst : label is "000006D000101000000000000000000541010101054545454545454545454545";
    attribute INIT_25 of inst : label is "68DCD946E4EBCF0EEE498C686B9D626F8619818080007C07C200984C15D40C10";
    attribute INIT_26 of inst : label is "CE57B18F66DF6733AF659FD96225DBD4722372CDB6B76E8CD18E6328DCECF9A2";
    attribute INIT_27 of inst : label is "D19B6EBD86716CDAE8E655BCB38B66D76732ADE59C7B376733AF619B76EDC35C";
    attribute INIT_28 of inst : label is "B374669CDB55BC3388E2CE04D76EDAE6F0CFBBA1B7EDC6CC732F1FC338F66E9C";
    attribute INIT_29 of inst : label is "EBE051D740A1E68046B76ECE655AC3E4F76A6CE675ECB5F1EDEE9CDB75EC79C5";
    attribute INIT_2A of inst : label is "02155A962587119ECB1A7DFF7F7053FEFE4F7CE792E0DB9B62EF3C59E78B3CF8";
    attribute INIT_2B of inst : label is "1111110000000011111111111111113FEC485111508D76FDB7B7567412048442";
    attribute INIT_2C of inst : label is "0A888CD41428888892222220BBBEFBEEEFBA22A0A28A288AA28A2288888A2B11";
    attribute INIT_2D of inst : label is "222222222222222202222222222222222222222222222231EBEFB6DBBEFB6A15";
    attribute INIT_2E of inst : label is "11004404404145B4151B051B451BBB19BB90546C146D146E2222200222222222";
    attribute INIT_2F of inst : label is "0820A2200080A0000088002D889D800001508A889D8004014000000040000000";
    attribute INIT_30 of inst : label is "A690A8150FFEA6ECEE8FFE3DFE00EF7275770770757EF936761231272F4D85D4";
    attribute INIT_31 of inst : label is "5545403E0ECEE3F3CEE0EAE4C0DC0888990DDC13CEEEAEE0EEEE8FFFF0EEAEE1";
    attribute INIT_32 of inst : label is "C007A62B0FCFFF6F1E2CEE2CE6ACEEEE0066600011660AAAAA4EEAEC3DFEE2F4";
    attribute INIT_33 of inst : label is "BEA7A435086CEEEEE8EE2AA2A2A9ABE7E0EEECEE6E88AA264466577737671990";
    attribute INIT_34 of inst : label is "000000002FFEE6ECEECFFF7FFF39EF7375775770FFFEF9BFFFDFFDFFFFCFFFFF";
    attribute INIT_35 of inst : label is "00000000000000000000000000000000C307723D515F71E033227941948A0284";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "087119CCD95EE30950E007001C0430100100100100104401C3C11036D3113000";
    attribute INIT_39 of inst : label is "7837C17CBF33C4BE7E666C978565DBE7913102004126CF024D9A01E00700C593";
    attribute INIT_3A of inst : label is "00180313F3E22357DF0920B2E067CF672DD9F92ECFE4000DE001ACB2F0017216";
    attribute INIT_3B of inst : label is "0031DD16492B724DFD3492E56FC955896040350F25601835879297C0A4430060";
    attribute INIT_3C of inst : label is "43C320E19070C878643D320120025FFFFF8122120121FFC09128102882809D16";
    attribute INIT_3D of inst : label is "402036EC0C4030C320E19070C87865E190FC320E19070C87A641D32C3B0C8786";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000A4D9B6F680E4811E03601E00FFC00086";
    attribute INIT_3F of inst : label is "3400000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "76D86BEB05E860CE1F522A83070E24550A04301982AAD4006E00000376D90420";
    attribute INIT_01 of inst : label is "81FF0195E676DA5152371FF70FE5CCE168373923EC70859AC6D93FC2E37D9F5B";
    attribute INIT_02 of inst : label is "491FCA366A93350E6EC22AA5365F6B2FB426997FAEDDCA9AEDC37E2946820D16";
    attribute INIT_03 of inst : label is "022F755F7FF55C44A011C9E72F536E674A34687EDA7B484AA003FDB44D909DDA";
    attribute INIT_04 of inst : label is "E1034E7C8C1796C7BEEDA6E8148B444428280508428AAD210050C6464671CA0A";
    attribute INIT_05 of inst : label is "03A91548883D107A241F112078D3022550051C0D21B3CDF5C8036957A9459117";
    attribute INIT_06 of inst : label is "CCD766BB354041260365CFCDCF3DC6767371BDBDC6F7B7583BB3BBC1DD9AAD96";
    attribute INIT_07 of inst : label is "F17C7610EA7C7610E26F8EC21E0A947E0FAA00043201F0AD0A1A95C25E01672A";
    attribute INIT_08 of inst : label is "A8AA1098001258AC247AF509F509E3D4FC2E52300E12D14214A9023FF156A338";
    attribute INIT_09 of inst : label is "D97201548D50607A1FC09339463D142C3A3A73A71D082A741AC2A8B025501DC6";
    attribute INIT_0A of inst : label is "2A6CDEF3DFFFB3692C748810089E95A01B2EAAEF07666AB45CFF7F97FCF30DF8";
    attribute INIT_0B of inst : label is "E16567518002003580D1ED5CD9BDF79FFF669799FEEEED60E942D851D2859677";
    attribute INIT_0C of inst : label is "DCB6B2E684400824A0CDFDD9DFFFB6D812811C3C747447C3F0FC40B6A4A0A40C";
    attribute INIT_0D of inst : label is "555DE6E35D5C573B90055C799BE6FE841A6FB6824B692926E7669FD5B1F96F96";
    attribute INIT_0E of inst : label is "0BA2BBBB0F31A26CC5E77EEF84DBA06EE5E4ADBB9FF9FF46A1B7292DCACD60A4";
    attribute INIT_0F of inst : label is "657DBB48ACDEF6DACB2BC4FAE948A4484E7EC57255634688C004E074722C805D";
    attribute INIT_10 of inst : label is "B48A400410D5009D4D4C1400C750036001495498B62136AB5FA43FB0C6AA84A0";
    attribute INIT_11 of inst : label is "090A8210854AA0825DC326192915505A12A5A92B08B00109692A000882038244";
    attribute INIT_12 of inst : label is "540835480F51177257C12990FBA0E8AA514CA441B15481090A8210854AA08201";
    attribute INIT_13 of inst : label is "BFB6F6C59B2A02F44BABAFC71C9740AA152D5C756805D4125444AD72F8711029";
    attribute INIT_14 of inst : label is "513D2F970CDFA95675792B1DBAFE4A3925D51410F31DBAFEA91E9A7B6292815B";
    attribute INIT_15 of inst : label is "81A00FC00712A1415534941022E5ED500070845CC02040AE76596FEDBC71F405";
    attribute INIT_16 of inst : label is "548DEFF7FD085856A8F05B6B1EB1D571FB60FA61E9B03711B5EA975E2C905F8F";
    attribute INIT_17 of inst : label is "9FED87FB73AFE2210A02120C10E3810FDB1122A14E09CA9744A8D04094485401";
    attribute INIT_18 of inst : label is "24895851A14A52C2E74E285EB7920CEF1CDADFD0286D821C7A5A9FB758A29020";
    attribute INIT_19 of inst : label is "68FFFD347FFEE15510976A869F0595E77B37DFB12140348802921029852A092D";
    attribute INIT_1A of inst : label is "0AD7A7A3314EC194DD888880CE9557F0478DC435886B7D110039309D13AC9FFA";
    attribute INIT_1B of inst : label is "C2CEB9BEF520223414A584B1E21131D0D12C0425285F4E614A14EF84220368C0";
    attribute INIT_1C of inst : label is "80A2B16C284428D4A6361C28C0659B2EB2EBB3F4180DDDDDDD997677766642AC";
    attribute INIT_1D of inst : label is "058CCF8892B5C8BB1BE374384443AC755ED4DB2ADA11712B61311E0A413D2186";
    attribute INIT_1E of inst : label is "D010A6A2286900023311800C35BADB5C341A1020914246A2A191E186F90F9217";
    attribute INIT_1F of inst : label is "30C0B75BB379A22951B50AD15285720252B0165ACFD2283F37E9DBA56DAA50BA";
    attribute INIT_20 of inst : label is "5A9154803009026125F0002910040484432000892DDB66E0B76CDF72376EDB37";
    attribute INIT_21 of inst : label is "9180F0100F002C13480303BF2420A80200080008459CA2C5E2E3FD6A7E202740";
    attribute INIT_22 of inst : label is "446840602102C70799EBBDF0312ED37C0800000070879010002508019CC10033";
    attribute INIT_23 of inst : label is "0000000001E0E0E0E0E1E1E1E0E1E1E1616060000160808F0E1603A09A103684";
    attribute INIT_24 of inst : label is "00000ED01000001FFFFFFFFFFFFFFFE000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "1696963440AB94A634A511554A1548BA8421E1008002AAAAA808000C15D44C00";
    attribute INIT_26 of inst : label is "B406A520342C95AC68C5248D12345033A320A0961A024178254B52C488CE904C";
    attribute INIT_27 of inst : label is "2D0495A904A4868592B5AD58A524342C95AD6AC52901A095AC68C12034128216";
    attribute INIT_28 of inst : label is "1A09C168248D08252DE294A82241242460925BD14168912A5AD2948252434128";
    attribute INIT_29 of inst : label is "824A0000949249280842412B5AD4822A424412B5AD48A964054178248D185290";
    attribute INIT_2A of inst : label is "0B9054200805ED059025563C1E090B54D5A6395D604892D25920102412048048";
    attribute INIT_2B of inst : label is "CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCABFBE0ABFEFFEFFEFFB24A1425011C65A2";
    attribute INIT_2C of inst : label is "AD55E56AAD755555599999A0B010010004033555D5D75D555447DF7457D759CC";
    attribute INIT_2D of inst : label is "99999999999999999999999999999999999999999999999FAAAEAABEAAEAB57A";
    attribute INIT_2E of inst : label is "FBE6A26A26AEABAABAA43AA47AA4FAE6AAAAEA90EA91EA93D999999999999999";
    attribute INIT_2F of inst : label is "0800222001E02000017DD55225AAF162FAAD1CAFAAF166ABC000002AAE1A69AE";
    attribute INIT_30 of inst : label is "40F0E97E09989198BB8BBA3DFE11899880880FF0B026603EEECEECAF2F4D85D4";
    attribute INIT_31 of inst : label is "F43541540B9981910770BBA1B2B82EEAFF0BBA13033330101010000000450DC1";
    attribute INIT_32 of inst : label is "FF5DAC40030111091A39AB1DF7BCFFFF11EE7BF2FBEF1776775763743DDCC0D4";
    attribute INIT_33 of inst : label is "FC06AC3F08311111107F6737F7ADEFE7E0777477321DD80D5DFEDCCC8CCD5DD0";
    attribute INIT_34 of inst : label is "000000002FFEF7FDFFCFFF7FFF39EFFBB9BB1FF0BEEEF9BFFFDFFDFFFFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000016BDC680989839508FEED06135CC3155";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "5211C088004FF0125AA01501128E1A38830830830A38401453C0FBD924881FF2";
    attribute INIT_39 of inst : label is "FC085BB49E000DDA3C062802DF790CEC8A70020D010A4F82149B03A915480D00";
    attribute INIT_3A of inst : label is "02691851E3E2222000200130A4A6C507C341F81A0FE0C9066C9067272648370C";
    attribute INIT_3B of inst : label is "AD33B85A6DBF5BE9F8A6DBEB4FD5812A22958022390ACAC5191C888321582B20";
    attribute INIT_3C of inst : label is "95924BC925E492F2497924FEDF6FF56AAD2801FFFEDB569400A264AD0AD2A460";
    attribute INIT_3D of inst : label is "423684CE094020920AC9256492B24949056924BC925E492F2495924922492B24";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000A149A5452174C10793B02A90203FE0F5";
    attribute INIT_3F of inst : label is "5200000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "56CA20F345AD56760F0ABAD96B0E1574B4CD90010A6992003500000FABA80044";
    attribute INIT_01 of inst : label is "8150419584E8F0AFAA6D17A146C1CAF478989FFD1D109D9B4B6BA4CBC7A4D951";
    attribute INIT_02 of inst : label is "025F587DD1DEE8A726A82AAF9ED5256A926AC8699659DAB2C969682242C30A2C";
    attribute INIT_03 of inst : label is "EAC86566BFE57558B21B41CD0E3D652542B081C139174A0261AE4272A3C70313";
    attribute INIT_04 of inst : label is "A17CC2ACF0C49255AC2D0653C5B1C38ABEEF050D088E48061167C1F351C54AC3";
    attribute INIT_05 of inst : label is "2A291948890112022481100400710210F41958A9A1220317E8402143D09EC43F";
    attribute INIT_06 of inst : label is "647323991D104134D2D307830613132322C4E8EB13A22C3311116198888C8B4D";
    attribute INIT_07 of inst : label is "E975F443E074F441E80E9E883C2B74B8050A02042041E02653909D215122D8E4";
    attribute INIT_08 of inst : label is "777000D34216787B847AFD01FC294FF0F42F63100C8044188610387D67C0E003";
    attribute INIT_09 of inst : label is "34C20D9487243E501EC32CC707FE288461B86BA11F0A0D589260B5B081383F14";
    attribute INIT_0A of inst : label is "0E24557A492499E51C1B081808DF641016182DA263323224B4249251266909BF";
    attribute INIT_0B of inst : label is "7D60E38534020419097531EC48AA93D24933B3EB9E6665FEE900BF15D2016B6A";
    attribute INIT_0C of inst : label is "CC1638E8D5606E920645556AE924924811215C2CCCEC8E58C2B08D9E7040AC11";
    attribute INIT_0D of inst : label is "59DC6625E946F738ACD22AF388E23B7956DBF8B6E3547CA2332F9F7D98E8BE8B";
    attribute INIT_0E of inst : label is "734CDA5CB76FCE4D6E7F6DF5D93FCC4D6E629ED68BE8BF0460932BAC4AD76D12";
    attribute INIT_0F of inst : label is "6164398FF8DCF639EEADD540FF15F8E7E675C78B89C1205DA041648C56272A9A";
    attribute INIT_10 of inst : label is "74B369D85179D2B15D59D5F49B56E745A547CB0A16A309116B8721182E494302";
    attribute INIT_11 of inst : label is "21424450914891177BC7363BB2BAFD1BDAD1BDAF09E2832CE94F7D2BD36955F6";
    attribute INIT_12 of inst : label is "6A2410DD1381802928DC9B45D29568E6C4DA1C2A818D81210244509148911721";
    attribute INIT_13 of inst : label is "47FF12530198C548A65E4B8A37520DCE2CC9C8D6D182EE2C747826515B0C5634";
    attribute INIT_14 of inst : label is "9A42709C8058004451C422004187DD1B0E46C1C7BA00418739687EA0EAD61949";
    attribute INIT_15 of inst : label is "9135910AEFA784CA6A720C0C3B8F04E3FF980E382AAD4A8C0026D1FFC06388CC";
    attribute INIT_16 of inst : label is "E36CB3D9EA25315C030410903E425D82D936412604955E14BF6AB65A2731B7DB";
    attribute INIT_17 of inst : label is "D2F794BDF94D0ABDC32B1D69BFC1D1FCCB545908CD0562109A12538E01B12160";
    attribute INIT_18 of inst : label is "06EF8AEEC46C20C35A670C5B131604455EDB55C198AD37F83AF3F9B21AD79163";
    attribute INIT_19 of inst : label is "F7CD587BE6D870B113F4B08584F585805E3BAF11A21C9A6AC1CCB6BCFF392837";
    attribute INIT_1A of inst : label is "08E2CAC471FF6484CB1BE1109DFEE8182F4FB0FBD9F7E93138283416825016B0";
    attribute INIT_1B of inst : label is "CAC891DD798D39D8D841879B4A8510A5E2F984A52CC831CC520407F0E8D3F69A";
    attribute INIT_1C of inst : label is "A853DDCC3667285025522F069A589EB8EB8E3178D348C8CC8C8A232223221C8C";
    attribute INIT_1D of inst : label is "F9E6C352D374D8E92F25E6B60243403112889184622CA091D13071855F0EAEB0";
    attribute INIT_1E of inst : label is "D501A7EAB3BE2B085C144107B49B8BF428FF1C068120111A35B178E6F9FF92FF";
    attribute INIT_1F of inst : label is "FB58174BA967BCB02CB23F0E2874B2A2F88F1158E99754CB7281C96FACFC2DB8";
    attribute INIT_20 of inst : label is "52911000070EAE0EC7AE0E2E3B1C84956A2A831805DB52E4176A59B2162EDA96";
    attribute INIT_21 of inst : label is "828CFE80CFE810D0200201980080B7E200B2A20C2A63AA03D013B7F5D646E040";
    attribute INIT_22 of inst : label is "503920006007C104910D0C60012E01AD087F800050000000003900010C500021";
    attribute INIT_23 of inst : label is "000000001D9D9D818100100C011C10101C0C10C0C00C4C4FE80E408A8E499392";
    attribute INIT_24 of inst : label is "0010166000000000088A80080008000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "5A0E0BA3B663FF13DB62C8A8F14CB2D7323E0C860001C71C7010000C95DC0C80";
    attribute INIT_26 of inst : label is "536558CDBBCED3976732D8AA7AA9DBA52AAA996AD6DABDB6BC87217676D4FB7B";
    attribute INIT_27 of inst : label is "B6D6FD1ECF59B779DE72ECE65BCDBBCED3976733DE6DDED3976733DDABDA6DCE";
    attribute INIT_28 of inst : label is "DDEF35A6B7C8A67BC563EB04FABDBE32D96ED2B2FB57E5A639768F6FBCDBBDF6";
    attribute INIT_29 of inst : label is "BAA851755030A2A0649BBDA72CCA65549ABB5A72CCA6565936BDA6B7C8A6ADE4";
    attribute INIT_2A of inst : label is "120E4FFF7FD3974FFF8FFF3C9EFDF5FE66EDFFE9BBB201C02F4D36E9B6DD36D2";
    attribute INIT_2B of inst : label is "666666777777776666666666666666FEAAFCFEEEFEE000000C930B655B0BC1B9";
    attribute INIT_2C of inst : label is "180A053FBBEAAAAABDDDDDEA1140540550141F7F5565D7FD74D55554555D7766";
    attribute INIT_2D of inst : label is "CCCCCCCCCCCCCCCCCEEEEEECCCCCCCCCCCCCCCCCCCCCCCDE505018240501A811";
    attribute INIT_2E of inst : label is "8C827427427EAA5BEBA6BBA6BBA60555557FAE9AEE9AEE9BCCCEEEECCCCCCCCC";
    attribute INIT_2F of inst : label is "088280088A4002222046644BAB2318C2123384212318CC9C80000009C90C30C8";
    attribute INIT_30 of inst : label is "C605AA81077EF770774664044411EE2471FF0FF0B895F818991111190D4F86E4";
    attribute INIT_31 of inst : label is "02D42839071767F78FF0F761F6FD3333330FFE118FFF3CF2F6F7B7D7F3FF2FE3";
    attribute INIT_32 of inst : label is "B054AED50E0FEE6F1E7DCD1BB330BFDD11CC59D0C8CD1776775763743FFCE2F4";
    attribute INIT_33 of inst : label is "014701750879EE6EE87F6EAEF7AD666760DDDCFF3E5DD80D5576667717667FF0";
    attribute INIT_34 of inst : label is "00000000277EF775774FFF777731EEEEFDFF1FF0BABFF99DDD9999999DCFFFFF";
    attribute INIT_35 of inst : label is "00000000000000000000000000000000183B46B44E4E91814C294F803B0FD7B4";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "1A11C0B4C04DF4007A2911003824A29A09229A29A29AAC144181FFEFF688150E";
    attribute INIT_39 of inst : label is "EE478B889F13E5C43E24148E584ABADEB16803650060C9D0C193822911003A90";
    attribute INIT_3A of inst : label is "0A050243E7E2237800000412343249C2E270D913C406881D68130966B409B311";
    attribute INIT_3B of inst : label is "819D9B4F249629A97D9249464BCC50A162503052A1281107215494A0250A2060";
    attribute INIT_3C of inst : label is "7DE73EF29F79CFBCA7DE73FFFFFDAADC0869037FFFFE043001502281A8121CA2";
    attribute INIT_3D of inst : label is "5A0605E6154031677FB3BF595FBCEEF2BF7657EF3BF595FBCEFD6536559CFACA";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000CC197FAACC74E83713F8320020000C95";
    attribute INIT_3F of inst : label is "9800000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "564A61C340A47446C25890095364B1201050120A04D22410F1020008669D00CC";
    attribute INIT_01 of inst : label is "125A4722757C589A2BB761274DC1CA64397CFDB30C3891CAD6596D892EADDB50";
    attribute INIT_02 of inst : label is "681802B5435BA1AA6CE02AA987740EBA06D2DC79A6DDC894C59B68294859083B";
    attribute INIT_03 of inst : label is "46502328332320CAB25518F46613273F02218B405C031029233A00B881C28281";
    attribute INIT_04 of inst : label is "04286A2CA08DB6C58F8E26C14191D0982241552C09AA45050B238545E7518641";
    attribute INIT_05 of inst : label is "8CA225110192036408D8204640172650C24E2CB5B6A412131068E0C069450032";
    attribute INIT_06 of inst : label is "EED7763BB4424CB44A8A2182203226666289B9BA26E628813BBB45099DDAAA28";
    attribute INIT_07 of inst : label is "C5616182C8E16182C8AC2C305889153141A86E4CA57A02A509D8C5AC5EF8B4A0";
    attribute INIT_08 of inst : label is "8AAA9B51265D338435A2892A8809062540A99B72521A110A0E903061230188A1";
    attribute INIT_09 of inst : label is "228A2651015223226D0987A5062420A083E00E203023AA41DB7AA201DE2A3446";
    attribute INIT_0A of inst : label is "256DEEC7FB6DB3C00090A3292A0217925451051426776AA1A2DBEDDED8032888";
    attribute INIT_0B of inst : label is "68B47515124A17660CF1149ADBD9FE36DB67801ADEEEEF038808E01F1016E766";
    attribute INIT_0C of inst : label is "F87EC8C04440000B85DEEEDD9B6DB6DB3B02105B77570F4D47D19C00ACA29C95";
    attribute INIT_0D of inst : label is "891DC6F1361CC63B8A0074E728CA3935627191326321F08EE6BFE2635EC26E36";
    attribute INIT_0E of inst : label is "596A0644264D8DDF7678ED1591220FDF7662848026E36C4065B64041F0C46031";
    attribute INIT_0F of inst : label is "CC8F190CAF0D77181D70C47F492650C48426152041894C88CC484864522CA24B";
    attribute INIT_10 of inst : label is "5BC18420444C0102020060128C807904121104BE7E24968C2802789096CB90A9";
    attribute INIT_11 of inst : label is "6DAEDAF3B6CBB632BB802401291405B96A7B9EA419C2830AB7848A110A892165";
    attribute INIT_12 of inst : label is "5028E1B1299191214310B65172A648EDB5B2A44CA1DB676DEEDAE3B68BB632C7";
    attribute INIT_13 of inst : label is "65B616F61DB04A11EC30668A204E0A8655A8888143DEDA52E4608452622D7625";
    attribute INIT_14 of inst : label is "CC83F0D9240FEB017C11A844B9015AF12C191410B444B90100E79D977C0A155B";
    attribute INIT_15 of inst : label is "A513CC98C7820DA839775819668165880002DD4108205088803A996D8577A6AE";
    attribute INIT_16 of inst : label is "9CC428944D2A511E01A1492061C608DBF370C17305B4CFD9B54A965A2572DF2F";
    attribute INIT_17 of inst : label is "66CDD9B36F1D0231C1E3189193859138ED162AA11E4B82420AA8920B9020140B";
    attribute INIT_18 of inst : label is "370F089085A2534A7C400E8A37123CCC1C5B1511998E3270B4A271DB389F92E6";
    attribute INIT_19 of inst : label is "FB8C467DC736F34732300934D4433E323BC1968D4052A0922290B248853861B3";
    attribute INIT_1A of inst : label is "2B56AC86361A0470000101328E154899688F00C70B8E99176869C4E19C30E08C";
    attribute INIT_1B of inst : label is "99249E0CB684B210C4A69513440D328284909C631D8075EDE6D38181A84B2289";
    attribute INIT_1C of inst : label is "8D836517A367B02024CBCA4209645861861870E1D129D9DD999A776676660AAB";
    attribute INIT_1D of inst : label is "41CE47408E73F9EC5B8B6234506820422945068214805102AA5E5AD849B424A4";
    attribute INIT_1E of inst : label is "E05286249128211AB2A08CB939B20914B0982084C12810140272E2E439D76C4C";
    attribute INIT_1F of inst : label is "B34A8180C362A04D19B022526295A40812147058D5C2EDC55A61DB04648B58B0";
    attribute INIT_20 of inst : label is "AA225109C3CC4C042430E7AC6409B6447C21161CA06D86F281B0D9BB01036C36";
    attribute INIT_21 of inst : label is "1E5EFEFDEFEE22489C04462736780000A80000A143D2AA2388489B2B6605340C";
    attribute INIT_22 of inst : label is "03440414418514032C4291060920180077800000287FB83806421C0230338046";
    attribute INIT_23 of inst : label is "002202021C9C9C9C9C1C0C001C0C0C10809C8C90809C000FE141040051012440";
    attribute INIT_24 of inst : label is "01010801010101000A0A000A00000000008000800282A28202220020A280A282";
    attribute INIT_25 of inst : label is "24949470C283A28210F6145448500921003FE0000003FFFFFD00FF1D15D40C01";
    attribute INIT_26 of inst : label is "A416A42240B50528C14436A82BA0915AAA20209828250A48414A528E185C0A84";
    attribute INIT_27 of inst : label is "4908230500C44816A0A51828862240B50528C1443912050528C1453240A08854";
    attribute INIT_28 of inst : label is "2050C258413878272DE09C8A450A09A1A29926C4248112085289C28862240A08";
    attribute INIT_29 of inst : label is "5B7068B6E0C16DC18A640A0A538688FA640C20A538688DA4C80A584138781393";
    attribute INIT_2A of inst : label is "2421544411056B56A21644C3E1B5A15541203A55488892925124922482449048";
    attribute INIT_2B of inst : label is "110011110011000011001100110011501000154504900000036D981645198494";
    attribute INIT_2C of inst : label is "1AA00695142000001000002AB400400500144080000000028B3AAAABAA8A2F00";
    attribute INIT_2D of inst : label is "0220022002200222202220000220022002200220022002315055440005546811";
    attribute INIT_2E of inst : label is "00085C85C85155515451C451C451553155555147114711460022020002200220";
    attribute INIT_2F of inst : label is "0DD55DD55C15555554000AA05000061500006150000614512EEEEED415FFFFC0";
    attribute INIT_30 of inst : label is "43EF015488088198BB0BB9BBBA11EF3CD9FF0FF4FEB5F838AA2EE66E2E4707F4";
    attribute INIT_31 of inst : label is "AC456BD50E8080808880C4C0C4CCEEE2EECEEE028CCC0CF0D4C484C4C0880983";
    attribute INIT_32 of inst : label is "150E54010F1101191C5DEE0EC9D49DCE22CC7BF242631BBAB39BAAA82AB02230";
    attribute INIT_33 of inst : label is "B402FBD508510111101919988088088888ABB8BB3E3BB80BBBFF7EFF9FFE6FF0";
    attribute INIT_34 of inst : label is "00000000AA2ABBB9FF4FFFFFFFB1FFFCDDFF1FF4FEBFF9BFFFBFFFFFBFCFFFFF";
    attribute INIT_35 of inst : label is "00000000000000000000000000000000B12BB904E54FAF41E42EF411941EE904";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "CA518960C95CE00974A225107D30E4C34C34C36CB6CBB5548041CD34931925A5";
    attribute INIT_39 of inst : label is "447FA18C0133D0C602622093A407A95F3D0983B481EBED83D7DB04A225103413";
    attribute INIT_3A of inst : label is "09124743FBE237D00000008272700DC6E579812B8C050A14B03300AA6818AB05";
    attribute INIT_3B of inst : label is "03026152492832480494928540091140CA60640E253032200F129100A60640E0";
    attribute INIT_3C of inst : label is "D392698834C41A724D3926D34D34D02A054D03269A6902A6818E050310381113";
    attribute INIT_3D of inst : label is "148EE4F50A04009069C834649A324C4834610688834649A324D390610241A724";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000BD7DA4443D6EC16602705A21BFFFFE20";
    attribute INIT_3F of inst : label is "A200000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "A490429A49A5A2DE4A69080B3F24D2101EC5BA0B5E9E7402740200025CD0048C";
    attribute INIT_01 of inst : label is "5BE908582562010C2BAD200209557F406225A49009268D3C9413297BC72900A6";
    attribute INIT_02 of inst : label is "446092B4591A2CDF6FC9D7E1855545AAA23BD54DF69DC084D3793864AA790B69";
    attribute INIT_03 of inst : label is "2ED23321021768C9E3555695559F6FFF26CD880990125884086053209176A8AB";
    attribute INIT_04 of inst : label is "43C45EFC91ADB6CCAC2D926B5DB766C8C8AD9BAC6DAAE76D9B66155555D3E659";
    attribute INIT_05 of inst : label is "5EA0750383534EA603A8F41D479376C5875A7EAA0556B612B32634C47B6D56A1";
    attribute INIT_06 of inst : label is "CA8654B2A15BECBE4A10559814D84CC44C1311304C44C12B33AA08599D519000";
    attribute INIT_07 of inst : label is "4BA1A0035421A0035C2434206969DDD2BBF96F5DA547407D2CB80781FE23A0A2";
    attribute INIT_08 of inst : label is "999E59F92F54019CB5D54A9E4AB58D2F28709B3B7E01D762DA3DAB4212BA556B";
    attribute INIT_09 of inst : label is "8017AF40395866E134ABBF050E536CD80B9789520A56514C946521DDA2A0404F";
    attribute INIT_0A of inst : label is "8448AA849249222DB118D7BD69AB1D9AD082040566754640816D36836B4D68C9";
    attribute INIT_0B of inst : label is "E4EC6D0F935A5CB01882109091552424924460957DBAAB0656010124AC0714FC";
    attribute INIT_0C of inst : label is "D0A4EA845C9F54042C8AAA9512492491B61764E8544458484290996496BA95BD";
    attribute INIT_0D of inst : label is "AB50945D7A89D4A16AD7786708822351164B74965B31E58444AEA003DEEB28A0";
    attribute INIT_0E of inst : label is "54496E2E6527E5555C55C8B9348225555C4E0962B0CA0D5A0925565494B54DB7";
    attribute INIT_0F of inst : label is "160C996B81085F3C38F09BFA0B182DA87FAC0C9676EDEDDA1482ECD138BEB322";
    attribute INIT_10 of inst : label is "728B5294DF5DDBEAB2B5A8B2CBA6F0AD97705CD0A4C1E06124024EB2995FA4E6";
    attribute INIT_11 of inst : label is "256648519349921EDDACA5652E63343B0AC3B0AD3B164958E56D100A8A08014C";
    attribute INIT_12 of inst : label is "80A68840904DCD61300A880CB59262C204404624958423256648419309921EA3";
    attribute INIT_13 of inst : label is "AE921DB00181918CA008D14F29CED9008954E4A089A4C488136A7EB9818033A4";
    attribute INIT_14 of inst : label is "0802F17845E09A838AC9AF4F03A17593D81CB514E74F03A18E2B39ACE40EB292";
    attribute INIT_15 of inst : label is "121311098986046D30D20408CA4D2C5007D1D92D78F1E3C6A82BABA482EBC48C";
    attribute INIT_16 of inst : label is "1CD470B858B08576DB933E0630634CE36A42014205B10365BF37F6D87984962B";
    attribute INIT_17 of inst : label is "20E528A9526B0E492997786C32894B28926992EDAE8DDF1958ED96DEB7759DD2";
    attribute INIT_18 of inst : label is "352C6B12ADD359DAE2D69C9E25B06AA9549C2E56020D865120065125D1123429";
    attribute INIT_19 of inst : label is "A28812514495A5FF76088CB6BC385421304105B36311FAD81FDAF26995E065A0";
    attribute INIT_1A of inst : label is "69FFB0AC37210F5930152B16AE4516B291AC758C29181153329D44A09414A024";
    attribute INIT_1B of inst : label is "2C02820827E4EA55A6B3B5FAD6128AAAAA08CE77985821C4C2E38994AE4EB3C9";
    attribute INIT_1C of inst : label is "BB8C0A1420F47B30D51604934946D41041041ED4F92DDDD9555577557755D994";
    attribute INIT_1D of inst : label is "CD6A1AE30E338A0D432942714D5837000800030010001C002B9092B8056C0297";
    attribute INIT_1E of inst : label is "B03AF44EB365666D85301C9CC12D5229B599618CC57D01B64384BAFC2FB524C4";
    attribute INIT_1F of inst : label is "AB5CE8340246E6ED5921645B62D5960722523552AFD641CD524452AD6913DAA6";
    attribute INIT_20 of inst : label is "FA075039C7282A8C3952EE5853D9972D46A0A2B53A000494E80090A869D00025";
    attribute INIT_21 of inst : label is "045E0025E0020000000000000004008AA4008AA26F82EE36952FFC486FACAC3E";
    attribute INIT_22 of inst : label is "00800808100A00FC0000408005B900007FFF8000000008080620000000200000";
    attribute INIT_23 of inst : label is "02202280A29E9E9E821E1E1202020212021E1E0E020282901000D00820000800";
    attribute INIT_24 of inst : label is "010100010101011FFFFD7FF575757FE08000008082A28280A28282A220200202";
    attribute INIT_25 of inst : label is "C8D8D86CDCB7E75664EC72D2CC168F4B7FC01FFFFFFFFFFFFC40008C1DD48C01";
    attribute INIT_26 of inst : label is "C5944732ED964630D95F328B622DB39CA2EE2D9E3B2EDC8B996C4B0D9B451935";
    attribute INIT_27 of inst : label is "917263656CC65DB2CCC61B2BC732ED964630D95F31976E4630D95E32EDC8B658";
    attribute INIT_28 of inst : label is "76E65C8B931B2B673FF59CD9CEDC98ACAF9976DB6CDB1C8B6319B2BC732EDCCB";
    attribute INIT_29 of inst : label is "4D38869A710D34E2192EDC8C61B2BE692EDDC8C61B2BE5C65E5C8B931B2B8399";
    attribute INIT_2A of inst : label is "0AA352CDB32671E1E6E16900808F2755EB7BBEE2D58CDB1B6092491249224925";
    attribute INIT_2B of inst : label is "000000001100110000000000000000FBAAA8EAFBBE800000012750B70B968762";
    attribute INIT_2C of inst : label is "580AAC55542AAAAAB0000020115555555556C080001000028B2AAAABAAAAAB00";
    attribute INIT_2D of inst : label is "0000000000000000020002200000000000000000000000100000100000012AB5";
    attribute INIT_2E of inst : label is "5555555555515555545144514451551155555145114511460000202000000000";
    attribute INIT_2F of inst : label is "080008800000000000000AA00000020000002000000204044000001415555555";
    attribute INIT_30 of inst : label is "A80000008F7FE6E8EE0DD9FBFE11CF3CFBFF0FF4FEB5F83DFC1DD55D180B8194";
    attribute INIT_31 of inst : label is "AAAA80000F97E7F78FF2F383F4FDDDC1FFCDDD17177738B0B3B3B383B3777743";
    attribute INIT_32 of inst : label is "AAA000000F1FEFFF3A31771FCBF4338B33883BBB8BFB1DDCD5DDC9DD58D5FFF0";
    attribute INIT_33 of inst : label is "AAA800000AFBEFEEE0FF7FFFF7AF7FFFD9CCCC444C22200999DD189B999B2AB0";
    attribute INIT_34 of inst : label is "00000000FF7FFFF9FF4FFFFFFFB1DFFCFFFF1FF4FEBFF9BFFFBFFFFFBFCFFFFF";
    attribute INIT_35 of inst : label is "00000000000000000000000000000000AA800000AAA00000AA800000AAA00000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "6F512DF2ED4DD6ED66A075026D30E4C34C34C34C34C3E66ECAED8D369A5DBE95";
    attribute INIT_39 of inst : label is "54F7DE8B81A7EF47034832D2F486897E6BCD072F8B369B066D320FA07502265B";
    attribute INIT_3A of inst : label is "000303B3E3F7FB50000000BA6066AA50E29C2514E1158064B80610AA6C02AB41";
    attribute INIT_3B of inst : label is "814001DA6DBD3BEA8696DBA7540D39E07670380AA5381C00055292A4A702E070";
    attribute INIT_3C of inst : label is "5318298D14E68A734539A2DA4DA4DFFFFFE08BA6D26DFFF045000181D81D9013";
    attribute INIT_3D of inst : label is "060795C46F098A9829CC14460A33050D1449A28CD14668A334539821A660A630";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000A6D3254C26C183EC0720EA07BFFFFE80";
    attribute INIT_3F of inst : label is "9200000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "76DB24C36CC94446994A3BD143429477A09D104D5A0C5000DE030004336D0101";
    attribute INIT_01 of inst : label is "80FF78F08056795D62239B7165C5C07628B5B24B0C98D18E4649AC89AD6D9B51";
    attribute INIT_02 of inst : label is "0056D9FC823E414C6D842AEDB4574A2BA4E3D97DA6DD9BB0CFCB782056826804";
    attribute INIT_03 of inst : label is "089A544D4A544514AE01C0C706716E0542B005ECDBF36802A0ADD9B63980080A";
    attribute INIT_04 of inst : label is "C840CC5E806DB6C5AEEF06F0C401618694E3FF0140020D01105440C0C0410000";
    attribute INIT_05 of inst : label is "2B049924A5214A429090148400E6001810010C1D03A207007249081441863104";
    attribute INIT_06 of inst : label is "666233119602801290515229128902222252AA890222253019992180CCC88944";
    attribute INIT_07 of inst : label is "2810100020101100293202200508BC4A0EA8020001C3002458880C905F20E426";
    attribute INIT_08 of inst : label is "888A004A4206C880000A25022509A091180651602C008000048B061AD4522810";
    attribute INIT_09 of inst : label is "945201924E91624046C0872102080028108A88A2460A28210A22808881000900";
    attribute INIT_0A of inst : label is "2A6C6446DB6DB14000169848020ED5D0028828A6022322251592490490200148";
    attribute INIT_0B of inst : label is "E0242404A40014200851450CD8CCB636DB62900DE6CCCCA22A12885C5420D31A";
    attribute INIT_0C of inst : label is "D91604DA9471C438C2C666588B6DB6DA1220520599998351545501B201202808";
    attribute INIT_0D of inst : label is "399C4233B4C4E6189E0016512ACABF3D02CF3C12C30C4182226396ED18F92F92";
    attribute INIT_0E of inst : label is "4769CC0C3600084445618E319804484445720DFF92F92C8321B6191846CE6000";
    attribute INIT_0F of inst : label is "3C318088FCCE67181870D64268006008C42D047F5CC3040C7C21C078B45D7F3B";
    attribute INIT_10 of inst : label is "F6B27BC844EC5210C8C90D141434A2412418C69B16A3690B5425FEB0FAC7FE82";
    attribute INIT_11 of inst : label is "4828929A246A24A3D532F19791999E7A9AA7A9A88060810DED0AEDBB90739816";
    attribute INIT_12 of inst : label is "3C2811DD2309D5715854BB10B1A4C0CECDD8B649819DB44868929A246A24A394";
    attribute INIT_13 of inst : label is "AE4916C9024980E152199F4506400082046C741072848C05C262BC328A384535";
    attribute INIT_14 of inst : label is "4242351FF44080C003BC021345A99A882C8074F37E1345A9945918646041015B";
    attribute INIT_15 of inst : label is "A1A50352818389EA51B51C17FB47BDC910EF87580E2C58A4002FEB924165FBFC";
    attribute INIT_16 of inst : label is "568462B15A05280400F7569050E5D567F364416505B81740B522C6183F90578B";
    attribute INIT_17 of inst : label is "92E584B9610F82253289083818A1818ADB5930800DE0820783AA500601B8607E";
    attribute INIT_18 of inst : label is "808C98604018108164699CCE3716066F1E5E7F20482F0314321315B61882F121";
    attribute INIT_19 of inst : label is "28AE751456CEC14D000C08039810F0C30F35D710A010A4280A83B4858227000C";
    attribute INIT_1A of inst : label is "0085A241B005E1D25C8388A00C2BF6B0920CC4108A213414401C3E1DC3BE1CEA";
    attribute INIT_1B of inst : label is "784619AEB4890C08302103F6EA011080801C142529C864694C10A88818946E52";
    attribute INIT_1C of inst : label is "8908925C402C0A108C0604AE52340288288203994A44CCC8C8C933333332008C";
    attribute INIT_1D of inst : label is "6186E302C1E0482B0BE1743707C80CFFEFFFFAFFDFFFD3FFBD717F90032C005C";
    attribute INIT_1E of inst : label is "D090A6292AA20E189FD1C40865B4DB1C18580C224108000A3410E0E038872464";
    attribute INIT_1F of inst : label is "2655B2593960E28954B2038618344A121821085CEEC36C463109DB06AD8A50B0";
    attribute INIT_20 of inst : label is "1A01900401100703ACE0020030042200C22025076C9272DDB24E582EB3649396";
    attribute INIT_21 of inst : label is "F9A1013A1013FF7FDFFFFFDFFFF00A0A8000A287C390C62052FADCBB6A406441";
    attribute INIT_22 of inst : label is "FF7FF7F7EFF5FF03FFFFBF7FFA46FFFF8808007FFFFFF7F7F9DFFFFFFFCFFFFF";
    attribute INIT_23 of inst : label is "88A8AA2A001C1C1C009C9C9C809C9C8C80808080808080800FFF2FF7DFFFF7FF";
    attribute INIT_24 of inst : label is "060E1FEE0E0E0E0AAAAAAAAAAAAAAAA8088888080AAAAAAA8AAAAA8A8A8A8888";
    attribute INIT_25 of inst : label is "320606004403B0A61EA000606B006890363FED8687FFFFFFFC04000C35F71F26";
    attribute INIT_26 of inst : label is "300134A00001918C0001A00040011A7B802882D100000320640310C00800C4C8";
    attribute INIT_27 of inst : label is "640C9000169400003231800034A00001918C0001A50001918C0001A000320006";
    attribute INIT_28 of inst : label is "00190320648000B4ACC0D2802003240000D000000000532018C000034A000320";
    attribute INIT_29 of inst : label is "0008000010000020000003231800000001003231800001140183206480007A50";
    attribute INIT_2A of inst : label is "3608016058518E63B0A33700809C50ABF5AAFBDD682A00C01C00008000100002";
    attribute INIT_2B of inst : label is "000000000000000000000000000000041500550114800000080100010817FA28";
    attribute INIT_2C of inst : label is "5AAAAC55542AAAAAB00000201555555555540080000000028A2AAAAAAAAAAB00";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000100000000000002AB5";
    attribute INIT_2E of inst : label is "5555555555515555545144514451551155555145114511460000000000000000";
    attribute INIT_2F of inst : label is "080008800000000000000AA00000020000002000000204000000001415555555";
    attribute INIT_30 of inst : label is "000000000111011155066062662202202222022022313035743FE66E2E4B83B4";
    attribute INIT_31 of inst : label is "000000000D9181130550D1C1D4644440664666268EEE6CF0E4C404C4C0880A83";
    attribute INIT_32 of inst : label is "00000000091101111C59DD1DCBFCB7CD11883BB989DB3BB8B33322646220AAA0";
    attribute INIT_33 of inst : label is "0000000008D9898991555444440444CFD9EFFD7F7CBB7C4733753EDDDFDF3AB0";
    attribute INIT_34 of inst : label is "00000000555DDDD9FF4777777733D66477771BB02237313FFFBFFFFFBFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "4800406C401B34000A201100010014004004004004004FFC0200725B6D800FFA";
    attribute INIT_39 of inst : label is "57904908011C248602386C0F284390AE092801648123C60A478C132019005D81";
    attribute INIT_3A of inst : label is "FFFD0101E3FA22AD55500420202285222740A03A050280294800A14494002234";
    attribute INIT_3B of inst : label is "843FFF2100091410830800A184020EA0201017D449084BFFE22081182101200F";
    attribute INIT_3C of inst : label is "2CD7166B8B35C59AE2CD712496DB300A0120004B6D93009000FFFE8028000FA0";
    attribute INIT_3D of inst : label is "EA0288C019007157166B8BB5C5DAE2EB8B9D7176B8BB5C5DAE2CD71D735C59AE";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000E478FBA7E43C052301C132000000017F";
    attribute INIT_3F of inst : label is "2E00000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "72492E492C92684B29944B6185932896C3261C4F5E187048D603000EAB2D0321";
    attribute INIT_01 of inst : label is "EDFF38F088766114422699312484C836289D1249E49AE08E42C8C49124448952";
    attribute INIT_02 of inst : label is "98964BDC8C2E464427842AED347D503EA9238F248248D9B05F91393263246985";
    attribute INIT_03 of inst : label is "D10AD88D5AD88624AF81484522222444932705B44B59389A218F68967C9C080C";
    attribute INIT_04 of inst : label is "9058C00AE2649274A4A5827EA0C269731533FFC166031833218840C0404C198E";
    attribute INIT_05 of inst : label is "2E2930498D031206B681B1B48CC6990E3DB3CF680D0154E8E4D9021400823C8D";
    attribute INIT_06 of inst : label is "4672339193369A132061D369D32993333274CCC9D333A63E119931F08CCCC9C7";
    attribute INIT_07 of inst : label is "31131206221313062B326260C70C1B4C4C04DBA210C1492A98800C1041012424";
    attribute INIT_08 of inst : label is "6661B6CC93824E6B63586C006C0119B03302756DBC24CC81A4C9C30A58542A1E";
    attribute INIT_09 of inst : label is "9870DB148C335A44D2761121319987031E9809808C8206060020068683080B30";
    attribute INIT_0A of inst : label is "322464424924997240139C9E8406741D038E30C7C33333261D000000063A8146";
    attribute INIT_0B of inst : label is "5B602034C9A124184859060C48C892124932908CE244469A6024869CC04D820A";
    attribute INIT_0C of inst : label is "4993A64D2771C43CF24644488924924CD049932C8898E36158D64092606C4240";
    attribute INIT_0D of inst : label is "10C84632D04432309709D8422A4A920A30C20B80C90701123267126610886486";
    attribute INIT_0E of inst : label is "8691CC0E120030444521843888047044452404EC864864A320920908424B30E8";
    attribute INIT_0F of inst : label is "3C21919870A52718187064822809A60B4829337FDC0202043E10827CA6595D34";
    attribute INIT_10 of inst : label is "729C294D64B66418484E0608601906F2499367899322E90D8439CDA0F086FF9A";
    attribute INIT_11 of inst : label is "9071230C492C48C1D512509290888A3C8B23C8B0C4790184E53045CCA0799802";
    attribute INIT_12 of inst : label is "7813125E470963409860CB2021488092CE5936910125989031230C492C48C1B8";
    attribute INIT_13 of inst : label is "6849E269034986A65269986186B06682344336135C80B435C24318248C388932";
    attribute INIT_14 of inst : label is "337C2113FCC088C003FF18374028A08880B76C5158374028DC6998A66071C949";
    attribute INIT_15 of inst : label is "CD4941648181126B919C27F7BB423A40001F7680864C990047C71A127B4D7B75";
    attribute INIT_16 of inst : label is "778442A152C524C50EF78E9180F86266D9283E38F89837419522D2493F901D0E";
    attribute INIT_17 of inst : label is "B64C8D9321279BAD1C9A11AC08A0808A4999359809E049B7F11A586609D0237E";
    attribute INIT_18 of inst : label is "E088C66C7348B4A1A4299CCE130606650ACEFF2848698114121114924E92F120";
    attribute INIT_19 of inst : label is "28A4D5145248001A880418E380D0F0832C24934CE10C1038C003992D6705D304";
    attribute INIT_1A of inst : label is "84816671ADC4B0D24C420C4809BFF5A09719C6398C736C1880162B19632F19AA";
    attribute INIT_1B of inst : label is "784701249DB24D8E116942648E210080806B21884347649B499C886F3B24E664";
    attribute INIT_1C of inst : label is "6810BA5C00241C3106260506643D238E38E3031F4C80888CCCC82232223274CC";
    attribute INIT_1D of inst : label is "248C4904F16C486D192329B737C04C0000000000000000001F506F801B080C5A";
    attribute INIT_1E of inst : label is "710083B3C4DB8E181FF1E7676495C9DE1E569E32018600CE199040A419132424";
    attribute INIT_1F of inst : label is "2E6512493B20DB3975939BB5CDA70E20D9ADCC4E6631888239108902C4EE7092";
    attribute INIT_20 of inst : label is "7293148F7D18DBFBECEDBA08DC73620446234DC74492765D124EC82E922493B2";
    attribute INIT_21 of inst : label is "0000000000000000000000000007FD5D75FDFD778490824862F80DB348736092";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000007F80007F80000000000000000000";
    attribute INIT_23 of inst : label is "2A0A08081E0202021E0202021E0202021E0202021E0202000000000000000000";
    attribute INIT_24 of inst : label is "000000000000000AAAAAAAAAAAAAAAA8088888888A2A2A2A2A2A2A2A2A2A2A2A";
    attribute INIT_25 of inst : label is "1206070634633C058BA088283B0C389E000000000007FFFFFC03FE2E35D40C40";
    attribute INIT_26 of inst : label is "33431DE9A760918E0C30EC0180060C2B80309873969A7126248320E0C600704B";
    attribute INIT_27 of inst : label is "24C49830C3BD34EC1231C1861DE9A760918E0C30EF4D38918E0C30E9A7126306";
    attribute INIT_28 of inst : label is "D389312624C1861DE45877843A7126061874D231DA4EF12618F41861DE9A7126";
    attribute INIT_29 of inst : label is "34D89A69B134D362649A71231C1863049A721231C186337D34F12624C1862EF4";
    attribute INIT_2A of inst : label is "551E0D7A5E918F2D3D2D2700006C52ABA1AAF398637A00C01F6DB6EDB6DDB6DB";
    attribute INIT_2B of inst : label is "1111111111111111111111111111111010045554448000000EDB026310155FFD";
    attribute INIT_2C of inst : label is "08000400002000001444446AB00000000002AA2AAAAAAAA82080000000000111";
    attribute INIT_2D of inst : label is "2222222222222222222222222222222222222222222222315555555155556010";
    attribute INIT_2E of inst : label is "0000000000000000010001000100000000000400040004022222222222222222";
    attribute INIT_2F of inst : label is "0AAAA22AAAAAAAAAAAAAA0088A88A8A8A88A8A8A88A8AD555555554140000000";
    attribute INIT_30 of inst : label is "000000000666477177066040442200111111111110000020202880080E4AC6A4";
    attribute INIT_31 of inst : label is "000000000E86E7D58EE0E242A0A8AA80888AAA268FFF7471F5FF3FF7F3FF5FD3";
    attribute INIT_32 of inst : label is "000000000E8EEE4E2C6A8A2AAAA8A6EE2244626040422EECA6EEE2EC6AE4CCC0";
    attribute INIT_33 of inst : label is "0000000000404444408888088088808A88ABB93B303B744EAAA822222A880880";
    attribute INIT_34 of inst : label is "000000005FFFFFFBFFCEEEEEEE228AB199DD9BB11115113BBBBBBBBBBFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "498076E6761918B60E293149119246496496496496490FFF627472592CE6DFF8";
    attribute INIT_39 of inst : label is "53B04871E0CC2439C198666A031B062C29160164092020124040262931484CCD";
    attribute INIT_3A of inst : label is "00071119E3E222A80000062D0100A02112082490411389231891E3019C482214";
    attribute INIT_3B of inst : label is "8C00030100018000834000300420CCE321319060119880003008C80233106200";
    attribute INIT_3C of inst : label is "2CF5967ACB3D659EB2CF596DB2492520A4720C4B6DB65239040003883880C0E9";
    attribute INIT_3D of inst : label is "0E328CC0931259F5967ACB3D659EB3FACB3F5967ACB3D659EB2CF59F71D659EB";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000E4047EE6E41209411082629200000000";
    attribute INIT_3F of inst : label is "1C00000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
