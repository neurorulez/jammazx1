-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "44A212715E5F7C71C1A49428B1054B47FF8451F4A891B426532EDB1795E00789";
    attribute INIT_01 of inst : label is "98AC7B4EA7EA9B7353567E0A86089A3C4A16806BC3C60C1E3C70F08FFF56B905";
    attribute INIT_02 of inst : label is "4C4F9D38C54569E720A366720953A9E74979BF4744000649CC51C54731471E05";
    attribute INIT_03 of inst : label is "24F8971479FDF3A4FB93D753CD045051C03B7BD3EE93EB9F652A7CFAFC9CBBD3";
    attribute INIT_04 of inst : label is "E59FFFAC880423AAF1AA6A147199CED4940E261977723FCDA38A4689874A9061";
    attribute INIT_05 of inst : label is "328A8194729DAE028402C006CFDECC55C43469761FB13A49B11D402229AF1073";
    attribute INIT_06 of inst : label is "1487D4211CB975E79195D54C0E8198A8D3EB9C5000B5002FCED22A1DDF276CAE";
    attribute INIT_07 of inst : label is "7F4D0AB4682DECC83790C13A11614C155ECBAFF3FCFB2F84C41E86A0092AC5AE";
    attribute INIT_08 of inst : label is "BC7870101C84D78859A0B9E8C9C85D91BB75497E8A2825DCCDC2DED193EFBA7A";
    attribute INIT_09 of inst : label is "BCF7ED90A8666633CC3D01F218B93AD806D86DAF34D3DCFD00EA8877BDF7C3EA";
    attribute INIT_0A of inst : label is "E7227EB11CF86B422234DE50E10C6215B3E15FD2148518914200BB23EAD2447C";
    attribute INIT_0B of inst : label is "2B4CACB0A1547BDFF40A2BA01737A2C79795B8BDB93D12B70BDBF51ABEAB5F9F";
    attribute INIT_0C of inst : label is "2AA2229F4D614543AD52D00022D25F216AA654A2A1D6D70D204050AD99D0F9FD";
    attribute INIT_0D of inst : label is "83BAAB28A077BD8053A061A9FA5A001114115D4C498A31112B5956CFFD987E6D";
    attribute INIT_0E of inst : label is "32A5FCE869703D095F7903FA2C45528A45EC1EC10816916FA57A7E444D78CC6A";
    attribute INIT_0F of inst : label is "C731CCDA5880FA27F4E96DFFE9730303135445F31355666BAEEC576B589DE57D";
    attribute INIT_10 of inst : label is "7DF71BCD296810128811023FB29CD6D9008055521578768F63BA55467E214FE2";
    attribute INIT_11 of inst : label is "36F9B9305DDABE33D9CFE064E41C0CBF4CC4735988EA713A98E6207C4A1A84B0";
    attribute INIT_12 of inst : label is "FD3F5959DEBA79DC4524F7E62703E3FE9383BC14CFFB8057EE8262DB78D3E69F";
    attribute INIT_13 of inst : label is "84010EEF9991FC7F23FA2944AFD6EEE94E9674FFC9AFFF5C2E27DFDFC48F32FF";
    attribute INIT_14 of inst : label is "D5A7621DDD34EAC3BBBF10024EF020187CDF99A3E055B390E88AC9C73963B20F";
    attribute INIT_15 of inst : label is "24C8200040E3B41FC90E235EB5758FDFB2A3F9F65F85FFF31FFF72E389008352";
    attribute INIT_16 of inst : label is "E6406000B080288419014801120151E001844280246400408042320800051830";
    attribute INIT_17 of inst : label is "000000000000000000000000000094E004231481442441410830000020440002";
    attribute INIT_18 of inst : label is "6F6D5D00003BFFFFFFFF1063FB4DD1794182D055AE31B4871452639620C7F6B5";
    attribute INIT_19 of inst : label is "88376B7577F73E022A23DDD7D7D7779CC2ED8E3A9C35F8DF558532A634074536";
    attribute INIT_1A of inst : label is "1750A0A0A0AC28290202E966D85996361642B8080016AD2AB5A01804C0626220";
    attribute INIT_1B of inst : label is "0000000228840500762951565454545548328CA1605A1A0A12828A5C5D931717";
    attribute INIT_1C of inst : label is "31115F5FBFDFDE92FE37FFB7DE973F9EAEA577A6AFF800060007FE07F8078000";
    attribute INIT_1D of inst : label is "24A70904AE3CC820046347290838045021C200A1E289199C0A1BAB6693754843";
    attribute INIT_1E of inst : label is "A9477CEFBA79DD15F457BB2B2964E48FFD59FB9CE7B0EC170808F7CF9FD06109";
    attribute INIT_1F of inst : label is "902546F6D6995CE591856337C5BFEC60CFECF4410F67F9C2DAFD18039DAA858A";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "B66727F2484910C3080026E47260A6880012301B76E7261022932C80221807A8";
    attribute INIT_01 of inst : label is "51C0FE507486738A7469401D5479D6025369CFB52A55AA52A5469E60007104B8";
    attribute INIT_02 of inst : label is "603604001889A3800D0E004C1A30204100402AA8885CA03028E3F2F8A38E448A";
    attribute INIT_03 of inst : label is "0A3B0C0D20242492920006CA1269C78EC00A1040A22AA0BEAF74820802002D75";
    attribute INIT_04 of inst : label is "DB212208BBB2EDB611DC06D8E692904A4DB8D752128CC80A10349F3209264E64";
    attribute INIT_05 of inst : label is "ECB45C1DB46210B0D65996F7E22801887668A313429AD01698D22B0500507B42";
    attribute INIT_06 of inst : label is "CADE66B6E000CE4B652FBE9352AA03114E14008F966869D65FA575A045473D58";
    attribute INIT_07 of inst : label is "83B1AF5A8FD140C9440A8A2363658C9613089900500823F2D98C1D92C11BD8A4";
    attribute INIT_08 of inst : label is "00AB33CCED19193592046103201AA5060C069688115116A04BCC04813DF130C4";
    attribute INIT_09 of inst : label is "FA8B2486458CA05190856C00DB43A32088A3B603896C6006983D1E87B40B1550";
    attribute INIT_0A of inst : label is "008D8806602323BBCC4B60CB64B99B5D468A82AD6F7EA3466C59B85AC50B398E";
    attribute INIT_0B of inst : label is "C4901125939994A0022EF4CDEA8134A60A5A21440A31A3541448A23952586065";
    attribute INIT_0C of inst : label is "44CCCB1C921F9A0A52EE2673CD88AEC69704ABCD052918D2B4EF6BB0002D13FC";
    attribute INIT_0D of inst : label is "CD485271C7B9454DE33DACB8C484DA2E60E2A435069427E6B4822A0319FC30A2";
    attribute INIT_0E of inst : label is "5F5A10039209C633A6361CD39D88A1148A71E30E3121268E49E4893E8A4D5994";
    attribute INIT_0F of inst : label is "108C214486F6D4CFC905800C12946A642DA9A66D65A980A2E515451D616E3E82";
    attribute INIT_10 of inst : label is "0005E090BCEAA24B9E8110A20C6450126909A77927ACA0C6905B68D80C6CC304";
    attribute INIT_11 of inst : label is "02202CBDE4111FBEDFD9D2AE2CB3509492994A25128D46A152945D4395A73B4B";
    attribute INIT_12 of inst : label is "80900405DDC48623985A24178668EC0063DFDEFB1802658C423D0D4593008044";
    attribute INIT_13 of inst : label is "B69762E20CB998AC05C86A9913B92AA9020AC908650BD4AD4A14966E22DF24AA";
    attribute INIT_14 of inst : label is "26000CE202491D144101324EE3295180050C80310B2020352B919F8B68A6A0DF";
    attribute INIT_15 of inst : label is "00009140800FDA711B28452006C0106003468A01805A0200A00600192523ED29";
    attribute INIT_16 of inst : label is "012390020C080028040000808902800062012035010140200410014432028400";
    attribute INIT_17 of inst : label is "00000000000000000000000010000A010314207C00023408618202004031A709";
    attribute INIT_18 of inst : label is "5FEC3D80002BFFFFFFFF310771F02DB008E480A7B033F1E80E710356620EE5AF";
    attribute INIT_19 of inst : label is "A2082A0A82A86BFD7FD7D7D57D57D78684BD9079A0F61E8CDAE62CC78200A417";
    attribute INIT_1A of inst : label is "81E41014101804060989303C8F0F33B3D3C31B0B0409B3E34DC04810C121E280";
    attribute INIT_1B of inst : label is "AC2AAABAA00080008040292C4ACACA4B82621206A988484860181C868725A1E1";
    attribute INIT_1C of inst : label is "582CE1144221555A30A02C08E3A18D47C672D953E3FD554E000FFF5FF80F8AAA";
    attribute INIT_1D of inst : label is "DB56FECE61ABB64A3E489095AF36A7EF35BF35DAAEDEC5AE777235516E1CE5EB";
    attribute INIT_1E of inst : label is "722D9F94D797637F9DA8C8FE72093B80002000238CE42AA6F3290C081069DAD6";
    attribute INIT_1F of inst : label is "274BD09B783268C7241F98DA62039B0D930332AEA98062B5800CF7FCF6755A7F";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "268B47F02222241042A024A261602247F80118C64CC35C0AF83C920630640784";
    attribute INIT_01 of inst : label is "48CC7F58B2E8BBC917092F0F9200FC747A48C424B93264C9972A5204051AA565";
    attribute INIT_02 of inst : label is "6000A9424CCDE22C682A0012B8180A22552814CCCC74A2CC2461ED6C9181778B";
    attribute INIT_03 of inst : label is "01109510080A959448B818512D404482E0108894548148B4EAB6C4123DB435AA";
    attribute INIT_04 of inst : label is "A7F7CF65001089CED30C021ED50E6582344EB40D6B56A56A87AFE7A8C3020241";
    attribute INIT_05 of inst : label is "8EA555ED391316809012A520A06745DEE65DE223C01AC21218430A8968489A71";
    attribute INIT_06 of inst : label is "43D134A4D42A7B7DB5BCF7D5542A0999C45280DD1CFE7B6C5037BEAC4B74554B";
    attribute INIT_07 of inst : label is "C0FD2BFAA169CEA961324B094549891464618BD4BD7187109002C0A401839004";
    attribute INIT_08 of inst : label is "B55E2199BB8F8FD8FA21388A129ADA45B536D62AD06A16D454260498B7FD32A6";
    attribute INIT_09 of inst : label is "068CA004012A6834D57A4A089271839C8CF2DF6FCDBE5414942F8AAFF0062B59";
    attribute INIT_0A of inst : label is "AFEAA7F544720ED1EA8DF0F3CB3553D5E552D15AD290B2B568120AF041501D7E";
    attribute INIT_0B of inst : label is "6EDBFBF772DDDE7226667E48FE113EF13C9F0B508B89B3F13532531E640B87B2";
    attribute INIT_0C of inst : label is "6FEE6FD2DD7CBD6C6D385C51EBF1B9F369B8B75EB6368D19CF31CCB087F553AB";
    attribute INIT_0D of inst : label is "E9E66FD166FDE4CCF884293B36CA8A2F562B78F9C737E2F5BB5E5A00D934CEA3";
    attribute INIT_0E of inst : label is "7B78B812DB69679BD7CF96F31958F336DB3DB7DB9825B4E96C96F166CBEFD9DE";
    attribute INIT_0F of inst : label is "5294A546DA343E6F2D85A41FFEB54D6F76DDE7373EDDC28D4DF81A5E7BB9F3DB";
    attribute INIT_10 of inst : label is "25EEA2452C42A4908C0251915E6118E349DD311AA1AC22C65052755002A8D8EA";
    attribute INIT_11 of inst : label is "44423D38EC033F946BD436EB28A85D8ADA4D29349A5F2793CA53E125AD694A52";
    attribute INIT_12 of inst : label is "5106D8DDFE26FA8FD50915C0815A08A091D5CEA91FF3C5954A2338CFD2910888";
    attribute INIT_13 of inst : label is "26815CFC01398462032803C03BB95555A306AD97656BCAE168525CBE643A1455";
    attribute INIT_14 of inst : label is "F3D076B81B6DCFD5790926CEB1D975397743A3CBC9250435D28C1FF40F614891";
    attribute INIT_15 of inst : label is "09000C2221037B1D1B0601FAD32DA8689BE0AB508F8AFAD0AF9510F60F79472B";
    attribute INIT_16 of inst : label is "0094084041700000C00410042020021C80588002820A82840124081080000108";
    attribute INIT_17 of inst : label is "000000000000000000000000020121001000810000418A9602442040948A0090";
    attribute INIT_18 of inst : label is "28F2C6000003FFFFFFFF900ECE60F38653AD15FBC9397BB49DBE1087201D88C9";
    attribute INIT_19 of inst : label is "90002A1006A02B006A022AD54002A9F56D0FC91F9239C3612589AB347A03CA67";
    attribute INIT_1A of inst : label is "2214000004040100C0C08A0381009070702061010480401C02005C0041746205";
    attribute INIT_1B of inst : label is "469101188000080800B031324D4DCCCC41926819665999999464630988A22202";
    attribute INIT_1C of inst : label is "784A3F5998CC18C90EB21318030398C8E231CEB15BFD082E000FFE0FF80FA440";
    attribute INIT_1D of inst : label is "D6F9BEB2C71685928F91A3CF734CA9FB676F45D10D1E8E19B583C2B34839EE2C";
    attribute INIT_1E of inst : label is "3AB42D0F9DC4C42AE5AF2C553A10FA07B900F40A10284A65CEE23031E3D9B7BC";
    attribute INIT_1F of inst : label is "05B89418E345600648ACD1474395A2C6A45A5675C64889270C55D19BE1ED2955";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "6240320B63C3A49A4AA2202D73E0226A8251100C4CE38462898C9B0611400780";
    attribute INIT_01 of inst : label is "9CF603BB37319CD3918B72CDA784CD939C8BE4998B060C583560DAC50510252C";
    attribute INIT_02 of inst : label is "12228906C44560A520220193AC5048724178166665E222584E7854FDB9E11A2F";
    attribute INIT_03 of inst : label is "0302C0CC8E8EBD52DC908C0B59014512C0001C90C48D481EC076F412109C1CE6";
    attribute INIT_04 of inst : label is "7FFB6BEDAB968DA240110CC5B398D412C9B2625B32526E54B2A2D98AA26A13A5";
    attribute INIT_05 of inst : label is "02191925B00D840034808C70002C4D56A164603610B00294B285080128115921";
    attribute INIT_06 of inst : label is "5D9BB1130D78232C9CD04ED6D6029888C869A2AD3DCE33684F96F728C26B4F1A";
    attribute INIT_07 of inst : label is "FEDBFF7C334CE5D7619AFB087164FCC7A65932F0AC5D6456CC07481002B75843";
    attribute INIT_08 of inst : label is "94B8F2A8BDADC4D8CCE510FB52481F82966EC0337C48070D47CE8471921B0EF2";
    attribute INIT_09 of inst : label is "C035E382046743A4553F23F859AEA8CBDE38DB2465B7CD58195DACBC55F5CACC";
    attribute INIT_0A of inst : label is "A52734937D19D0556665BE55E14CD7587166C5AF7BDEBAF74E83801806400CD8";
    attribute INIT_0B of inst : label is "665D8D923AC4731BAAB7670ECF3477756FFB3C5DA72FF76745DF5378808A1597";
    attribute INIT_0C of inst : label is "722364A65F2EF92C4F1C95DD6656B9627898A77C9627C77AD6BDEF79A53979FD";
    attribute INIT_0D of inst : label is "2F3209857EE7320DDAAC095562D3ABEB327C4B5E5B97E2B3A3CB0E518B9D5861";
    attribute INIT_0E of inst : label is "7760CE50CB2B7159194BD73755EAB5538B8DBCBBD97CB7F32EB2F3FEE329CAD6";
    attribute INIT_0F of inst : label is "5294A5C2CAB0B36065D7ED1E98B9C3F212C4599212C4760B4C8A165EF5BA62D1";
    attribute INIT_10 of inst : label is "35BA32E524602424CC09403B927018620F8CD51805F97446000B440E86C8A988";
    attribute INIT_11 of inst : label is "4C409D03DC977F61A10532C1A2A85A8A5CD47B59A8E37938DAE6207694AD294A";
    attribute INIT_12 of inst : label is "53024E4E72C2C8A8CD433976B66206A0B850606C4859D5B5418CD1C2D1B10988";
    attribute INIT_13 of inst : label is "2B3605054D968D874D7CE8151DF47FF8E58465D5E6A56A7C68574C9F600FB855";
    attribute INIT_14 of inst : label is "B145C6357165BD91892BAF6C159D6C185C4A618369B5B59879BB0DC6454FF040";
    attribute INIT_15 of inst : label is "3020001450C3EB3BCD66A64C912488C83F61BD9528F28E9508D23453D6BD56AC";
    attribute INIT_16 of inst : label is "4240450830027080100166024000018008045B4810042048008A002800A00093";
    attribute INIT_17 of inst : label is "00000000000000000000000000008412002800FC681401400000002000404800";
    attribute INIT_18 of inst : label is "086905004023FFFFFFFF00C2C049A0E021854883852177A28D70500E01858695";
    attribute INIT_19 of inst : label is "7AAA84BAA84A81AA84A8006EEEE8018C054D05198A30F0330180520488069403";
    attribute INIT_1A of inst : label is "220448484040101244C400218908327252088202000000000000000040036CAE";
    attribute INIT_1B of inst : label is "EC7BEFB0000002020000212048C84848010A4010643919190C44408888426242";
    attribute INIT_1C of inst : label is "3047116DD2E9AF5C285B5ED8A1CEFCFF5B9F9D9E7FFD5D7F555FFF5FFA8F9EFB";
    attribute INIT_1D of inst : label is "DCE912E79E9C3799898D9FE6B5C8DA95C644E44FE5126E7B19E55EBB23B9DEEC";
    attribute INIT_1E of inst : label is "5620819FC990E6A2788FBC45D601398AC68800808220121BA7845A34E9FCAF5B";
    attribute INIT_1F of inst : label is "33AE9428A112A00407A84FC743D0195D1179167F9F602F9B2D45A75E416D3925";
    attribute INIT_20 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_21 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_22 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_23 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_24 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_25 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_26 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_27 of inst : label is "F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "E8CC70027C7DB2C308C28B446B62B42AA95BA859767C4B5822B80009A8280781";
    attribute INIT_01 of inst : label is "0DCE8058526702C92B28265DE385DCB6592AEC108952240814205244A52B84F9";
    attribute INIT_02 of inst : label is "12B68805EEEFE9B081482080862240D2045954CCCE63530126EA4D6C1BAE064B";
    attribute INIT_03 of inst : label is "4F11D9DCB0B6E916B4C2595A0200018AC020B481942D40D4D0B6671011BCB5AD";
    attribute INIT_04 of inst : label is "48009209001289B40D2C0E4C91D1948854963050D0983A4E9882458A8B245A56";
    attribute INIT_05 of inst : label is "44901A41B462C02072495EFD96795FFFC18EE93F88F9140EF9122A15907819C4";
    attribute INIT_06 of inst : label is "4A1EC2140C99636DBDB516C407207DDDDA419B9C302CA5764D36360BDB651072";
    attribute INIT_07 of inst : label is "C1196B70ACE18C8B763A4BB0664CA9921B4D90B2A9592692890CD2B007911C26";
    attribute INIT_08 of inst : label is "B440673339EDCDDAD809B200C35C4A94E5E6C8A059E2070C9815988B021E2056";
    attribute INIT_09 of inst : label is "428B7934654DA6D7049A4E1A9155819BACB8636C64C60CA05C0D9028580AB559";
    attribute INIT_0A of inst : label is "3163A5B10CE980556224B001C404574D6552C1085290B0810C49C81D465B6C50";
    attribute INIT_0B of inst : label is "684B1B3066CCD6345324662CCCF336E2AC5B16579B11BB72E5045B3910D4C54C";
    attribute INIT_0C of inst : label is "3667759C4ACA3CEE6235C91462C6B67B11F8B01E77310CB4A52108B790304FA8";
    attribute INIT_0D of inst : label is "2D6623897EED66DFD1152B33C2792C8B1689191AEB5608B128B27B4B1136F169";
    attribute INIT_0E of inst : label is "2362B652C9CD63594333F667198CB916AB1BB5BB5BA1B00E26E2408ECB7980D6";
    attribute INIT_0F of inst : label is "084210F2727C5760C4859C909CAB8932B2CCF332B2CCCE66259E4D0085B4C2D1";
    attribute INIT_10 of inst : label is "27266DB494B203495C0D3826D4683BA32D8D227F838C1CC74143134A5CAB9B29";
    attribute INIT_11 of inst : label is "12423A229D6DDFD5683732D1D92F58AA4A4D213098572B9588436028C7318E62";
    attribute INIT_12 of inst : label is "5402DADA23424AC8460E6D5DDC6100AB4D11280D82535FCD4BFDCFD2F0C90A48";
    attribute INIT_13 of inst : label is "67353B9BBD71990D28DEB717A03DD555EB9AC495751BCA796012599056CAA155";
    attribute INIT_14 of inst : label is "B3FC161B0364CDD50909AFDD1E597B259344D26C4D201E08523185F56FA952B1";
    attribute INIT_15 of inst : label is "0400D18000008410046882DDB36D8C6CF3603BE22AA2A8E22A97F39D4631672D";
    attribute INIT_16 of inst : label is "802322000608804100C088000404100024830410643041202800514054029600";
    attribute INIT_17 of inst : label is "000000000000000000000000600008440301000103222409D0A201000A113001";
    attribute INIT_18 of inst : label is "536E2D80003BFFFFFFFF61E918910C061C408405B49AB44A424E4B76C3D2374E";
    attribute INIT_19 of inst : label is "0400000100000010000000001110018B80ACD4D829B60E8CD83684D912042654";
    attribute INIT_1A of inst : label is "42004444444311108404062008085212320A430304000000001FFFFFBFF87000";
    attribute INIT_1B of inst : label is "56D54550011A000000102120C9C9C84811064310A40929090048408888220262";
    attribute INIT_1C of inst : label is "1A0BE736D74FB76C206CCD4AA39CE6F5F9FCFBD963FD88AE222FFE0FFFDFF551";
    attribute INIT_1D of inst : label is "C4ED12339A2491058914ADEE7BE9DC93E644E4544D12A64F3D9EDC9940889F24";
    attribute INIT_1E of inst : label is "B034ED29704496EA65AD9ED530097A8AD518A78A14C8021FF7F809A4C9DDA379";
    attribute INIT_1F of inst : label is "273C90D9E34468D20A0F964C036D90069DA2D374DB25B42927B4D399E3EDBD55";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_23 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "AC66268B8484CAAAAB601B654BE6B6AF4DDBB9E147C8008106B36D9D2D37FF81";
    attribute INIT_01 of inst : label is "45CA86D5605436A0BAAC04DD413DD626D5A8ED900040A0428008025A9BB994A8";
    attribute INIT_02 of inst : label is "B81B92720889B4CA4DEA0700E93313449A42ABBAA9720491A2EA296A8BA8142A";
    attribute INIT_03 of inst : label is "08D1CCCA1213225293237D4A8065B2CBFFD4D32699329194A234886469253DE4";
    attribute INIT_04 of inst : label is "490410093B5267C1010D2E4986949A0A4494D8D04E24C999151485332D265A97";
    attribute INIT_05 of inst : label is "3492484CF81289127249B4B281A8A0890B28B4D303980E01980A29355A4E190A";
    attribute INIT_06 of inst : label is "4A480212400862698D9086880EB1411160880AAC512AB54DB900B414676FBC46";
    attribute INIT_07 of inst : label is "3E112B5040C1CD9B6A364B51234488B24892900160E24A128890CA924995895D";
    attribute INIT_08 of inst : label is "2980E31329290952930428C100818203250E80409A412F4006958180B0106020";
    attribute INIT_09 of inst : label is "7A482322448260B488B227E851519113ADA2824AC90440008C8D184841F71351";
    attribute INIT_0A of inst : label is "4A6EC9B7202350156E400ED54541D74B46968A4A4294A1022449B91BC48929A2";
    attribute INIT_0B of inst : label is "449110294A8894200AA57444E80174AA693AC4200A53A7484224A23C01000824";
    attribute INIT_0C of inst : label is "44445534924A084B422481146E96A04A1126A10424A10814852908B4022090A9";
    attribute INIT_0D of inst : label is "654442974AA94D4CB914EBFF549128CB764613509A5408B7D09228047B15D422";
    attribute INIT_0E of inst : label is "43410290124942518242545358AAADD0AA17A53A5120020A48A484969A5D1A94";
    attribute INIT_0F of inst : label is "00000064925554404915A02510439100808CE320808CD0121518A484052482FA";
    attribute INIT_10 of inst : label is "C947648894EA136DDD9BD2226460BE8B29ACA33993ADB1E628612048206AB906";
    attribute INIT_11 of inst : label is "20C37A62AE510132F8294EA3527255D49209082412040A0100004C04A4210A52";
    attribute INIT_12 of inst : label is "F01C9493BAC499181B01A69292C0ED710B93BCD859E3D587462D1BC28B070C38";
    attribute INIT_13 of inst : label is "AB9321017FBB4884044C6A4813B91113A306292E753814A80D70952AA25AA0AF";
    attribute INIT_14 of inst : label is "B31C02A501292D8318156ECE30255146A5849424892FE1BC11901A54AC66405F";
    attribute INIT_15 of inst : label is "C9800840052E906DDF246C9122493171874ECA20310113201136109114A45489";
    attribute INIT_16 of inst : label is "0C90980200A10112AA22000112D1220040088022008982810044080000002844";
    attribute INIT_17 of inst : label is "000000000000000000000000000300002004037C80899A920010308004220082";
    attribute INIT_18 of inst : label is "807006FFBFD7FFFFFFFFEFF00C02020082102201C044381021808407DFE00801";
    attribute INIT_19 of inst : label is "02200802008A88200800000A0A0AABC0100E201C403801002008010041F81888";
    attribute INIT_1A of inst : label is "00000000000000008080020081803030702011010000000000000000000060A8";
    attribute INIT_1B of inst : label is "451111100000008008020300414140C000020200A00808080008010100000000";
    attribute INIT_1C of inst : label is "193C02926134924E5420200F7755A8D1EAF5C89A83FA080E888FFE8FFA0F8444";
    attribute INIT_1D of inst : label is "FA5497D3496ADE3B4E38F5AD6BA5F4AB8525A57AA297C5223A1AA511FE0CA422";
    attribute INIT_1E of inst : label is "39C78DD0827F5AB545D40D6AB96FFF8F21593F9FFD748207FFE00103070C52B5";
    attribute INIT_1F of inst : label is "E085FA1FD7BB7508FD143AF8A501DD28D0070950010202F046025A91AF8E31EE";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_23 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "011082882222261864A2691039321067FBC884C00257FF7EF92A49040128079C";
    attribute INIT_01 of inst : label is "9CA6041B0731A0D38982724D86449D101C81E62DBB366CDBB36EDB25FF814206";
    attribute INIT_02 of inst : label is "3106C942444571A53220911682880A62546896666476124C4E5824ED3963F68B";
    attribute INIT_03 of inst : label is "111C61240808B518D898C8A3599A08A0C0329A94D48948AAFAF6C6F23C9435A4";
    attribute INIT_04 of inst : label is "25924B2FC41911BEF990D104B99CC4630A13371B68732D42C3C6C9CC9291A071";
    attribute INIT_05 of inst : label is "474B616A37EBAE41092462109A0D6445830471B2049032329033841028C17C71";
    attribute INIT_06 of inst : label is "636138C924486B6D99B6DEF42604C888E264888E300C617B7AB6F66D6B6308C2";
    attribute INIT_07 of inst : label is "C2DCE771AC5DA4C76192EB0D9CFA9F0D65454251A77514D9E603614D8140E620";
    attribute INIT_08 of inst : label is "BE3A78001585C59859383DCEC08BB509B326C1B2DBDE07647D445C1F921F13E6";
    attribute INIT_09 of inst : label is "01ACA1A91237C860F6759A093C62C8D89C30DB6ECDB72436A23DC1BC040D1ECD";
    attribute INIT_0A of inst : label is "2732B5B994190241732DB071F32E42707160E52B5AD6BCB9B3248C0950F6CE7B";
    attribute INIT_0B of inst : label is "72DD8DBD22C4731762347752EF9136E30C9B0C9C8B19B36149B3599BFEFFDC96";
    attribute INIT_0C of inst : label is "72232C86DB616B605B13301072F2BB62D8B02CB5B02DC6F2B4AD6B7C89B36557";
    attribute INIT_0D of inst : label is "53335B5162E73C2EB5C2601176E70C0B9B1AC8D8431620B916D98684F1AC5E33";
    attribute INIT_0E of inst : label is "6F66DE40DB67718ABBDBB7620E08B1120B8CBC8B0EA5BD736EB6DECAC36DD0D7";
    attribute INIT_0F of inst : label is "42108466D90073386DC7E473D9338B2212C461B212C462191C8832C630B25AFB";
    attribute INIT_10 of inst : label is "3DF6D6D6622069244A09083B576C1AD1858E38D1495E504680DCADA433208DF2";
    attribute INIT_11 of inst : label is "CF44BA08AEC761944B15B2FB68295ACADEC77B1D8EE379BCDEF63376B5AD694B";
    attribute INIT_12 of inst : label is "7B0EDCD932D6FCE8E51135F0F00613FD9901292A0FFB03BD52050160F4BD11C8";
    attribute INIT_13 of inst : label is "00C94D8D0C18EE76136D20624F7B2AA8A50D6DFFD2F66A6470975995ED95BA55";
    attribute INIT_14 of inst : label is "B1A276329B6D9DCD383EE36FB9D17008F8779097E495E81D2C4C0A4E07D2A101";
    attribute INIT_15 of inst : label is "000100073072529E0E9732DDB16DCFFF937379B06F84FDB06FFA50C70420440C";
    attribute INIT_16 of inst : label is "1240000418000C2000094204C000082018147240020000480438008FA0F54002";
    attribute INIT_17 of inst : label is "00000000000000000000000008041623C0884080500441400200000000408410";
    attribute INIT_18 of inst : label is "7F6FFD00402BFFFFFFFF100FF3FDFDFF7DEFDDFFBFBBB7EFDE7F7BF6201FE7FE";
    attribute INIT_19 of inst : label is "AAA00AAA00AA8AA00AAA0000AA0001BFEFEDDFFBBFF7FCFF9FE7FCFF3E07F777";
    attribute INIT_1A of inst : label is "40000808000200000080040001005010500141010000000000005C15C17060AA";
    attribute INIT_1B of inst : label is "44514510011020000000010040C040C0000A0000202828080800010100404040";
    attribute INIT_1C of inst : label is "3008BE590880596CDE3797BA293631196CD626DF5FF8080E000FFE2FF88F9451";
    attribute INIT_1D of inst : label is "C1F2561F2CB924D36ED3A614A592B2A79C95B7D384DE9DBEDD6BB237497BFCE3";
    attribute INIT_1E of inst : label is "D80830A6CD1479AA98A64D545890FA8FFD20F50A568801F803FFFFDBB73C8E52";
    attribute INIT_1F of inst : label is "12C614285D45A8F14982D30341B62AD126CA659B2D82DBA29AD924579096D654";
    attribute INIT_20 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_21 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_22 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_23 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_24 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_25 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_26 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_27 of inst : label is "8888888888888888888888888888888888888888888888888888888888888888";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "420100802222A41040E8000011400247FB8010C2024000000128000D08000788";
    attribute INIT_01 of inst : label is "D8A4744A3720A25B1903720CD70089104803C009B3664C9B3664CA05FF110004";
    attribute INIT_02 of inst : label is "2102AB02666770AD606001369A101822C4289444447402D86C51A4E5B1415299";
    attribute INIT_03 of inst : label is "00180344888A911048B0D1C159002000C01688B04589586A4A7256F63C941084";
    attribute INIT_04 of inst : label is "2592CB668010018004BC0204318854420C32320B6A76244887825C8883020023";
    attribute INIT_05 of inst : label is "038B4368300BAE002000A85001456664C28670B2009016109013100078417831";
    attribute INIT_06 of inst : label is "4343108164482924B8A65E541602CCCCE16480981024232D3292722D6A271C42";
    attribute INIT_07 of inst : label is "424CA730A45CE44F2190E90D15AA9515254586D1AD7516D14407838000004014";
    attribute INIT_08 of inst : label is "9C121000348CC488C928188AC082B501B32640B6515A06641544E89287CC22A2";
    attribute INIT_09 of inst : label is "002DB0802003683054250008286708C89890492484932412C01C88B3B40713CC";
    attribute INIT_0A of inst : label is "2F223491141900C122249010A10C42513162452B5A529891A290820820C00472";
    attribute INIT_0B of inst : label is "364C8C9D2244731322345362A59032430599181C8119932381935B1800003CB2";
    attribute INIT_0C of inst : label is "22236C924B612B605B13B01022509122D8B02C95B02DC6D2B5A529FC89917055";
    attribute INIT_0D of inst : label is "4333595122673CBAA5804022327608091C0AC9484912009116D90685E8A88E31";
    attribute INIT_0E of inst : label is "2722CE404967319EB949933204089116098D9C891AA4957926925E4A4934B053";
    attribute INIT_0F of inst : label is "421084625800736F24C7E477C8318326364461963644720B0C88164211924A79";
    attribute INIT_10 of inst : label is "3DF2D6550061000088090019134C1AC115083153017C70860048ACC4360114E2";
    attribute INIT_11 of inst : label is "0C409A28AEC6608402F4B24A082BCACA4EC67B1DCCE371B8DCF6227294A5294A";
    attribute INIT_12 of inst : label is "7B0E4C4844C27888470015F0704003FDB840420007F901314205016050B50188";
    attribute INIT_13 of inst : label is "4480E66634096452022C24405CD92AA9362624FFD3BD2ACC200748B1E0151A55";
    attribute INIT_14 of inst : label is "91A6621399249CC53C3FE378A8D332187D7781B2E49F200FA800020A0862A020";
    attribute INIT_15 of inst : label is "066294004260EF0F0612224C91248FFF9323F9900F80FF902FFD50C204204408";
    attribute INIT_16 of inst : label is "01200558060AA201408020000828000220610815952441303301106011000210";
    attribute INIT_17 of inst : label is "000000000000000000000000000000001000807D0402042D2C82C04013140068";
    attribute INIT_18 of inst : label is "00E000000007FFFFFFFF00000000040004000001800030000100000600000001";
    attribute INIT_19 of inst : label is "2AA00A00AA0A8A0AA0AA000000AAAB80000C0018003002004010020080000000";
    attribute INIT_1A of inst : label is "000808080800020080000201808030703000000001000000001FA3EA3E8FEA00";
    attribute INIT_1B of inst : label is "1404005000050020550405014141C140200A0000202808280800000000404000";
    attribute INIT_1C of inst : label is "3008BE4B0180CB68CE1793B26A72130BA46266560FF8A2AE222FFE0FF82FC100";
    attribute INIT_1D of inst : label is "91F6549E2CB984D26ED32235AD32A6A535951F13805C98B0503992264163FCE1";
    attribute INIT_1E of inst : label is "681C1682C8547B001C06CD00E800F28FFD20F50A562003E7FFE003DBB7380E52";
    attribute INIT_1F of inst : label is "10C6A4301E01C0010986D10101B2880382CA248B6D825BA69AC9305710926340";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_23 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
