-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity rom_cpu2 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of rom_cpu2 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "96F616B3B52B61651A7E46424E4671712C4B0DDD63F6EAA56D2DFF5B5D243758";
    attribute INIT_01 of inst : label is "F4F0A3C2D4A2C2799F5850C9C73E598F707389CA396712E2C5CF042595E5BD87";
    attribute INIT_02 of inst : label is "AA5D78FD5A146157924FF24E213F5E54A15613B656E251BD3B9E4FF9CFCF1934";
    attribute INIT_03 of inst : label is "4BF947073A4928251552951498F362A763EAD7FD27957652FF2555C71479A6B3";
    attribute INIT_04 of inst : label is "6925A15954555ADC5940857A2E8959491C1CC9473CA7552E5470735492864E8D";
    attribute INIT_05 of inst : label is "B727AC4A1284A26D656D656D3E43D73D63D53D58FAA6996956956956956D5859";
    attribute INIT_06 of inst : label is "CB0FB185CF0817F97FB95CFFFFD9F2C9C89C28273C20561CF0A1865A8E81559C";
    attribute INIT_07 of inst : label is "05E4D20E4EE711B74585CF0815A4D2C0A173B8254A4A425155D512C4B12D49C6";
    attribute INIT_08 of inst : label is "D3CC4BD49A7D994B460A94602C9A5AC99F99352E8250C6268294BFFF19054B2E";
    attribute INIT_09 of inst : label is "F468AEAA68AEA25635A2F5A2E529293B5C2111676492D7F97E36A464246424A7";
    attribute INIT_0A of inst : label is "5575D69EA6D98796E4B96E6B9AE4A12B385A9B9F4E7A2AA52974DF245125B4B3";
    attribute INIT_0B of inst : label is "AD8FF7BE5D2415E9550D90575B5263402636236A42555A4237D5A423795A4237";
    attribute INIT_0C of inst : label is "50541FE2A107A07FDBD91D41575A5553929298D64A9B42D694B85D43E496DCE7";
    attribute INIT_0D of inst : label is "0267DC6541E69898C9A98E4B566376401001CCD8894450018896BD01FF6DED47";
    attribute INIT_0E of inst : label is "208D67AAE4209900005115649FD29F6712F9D2E2A6635DE1BD8D8D29C2026502";
    attribute INIT_0F of inst : label is "D7D279C8D9DC714456965925276492DC8D2B92D4A082359EE96768DC4AE4B528";
    attribute INIT_10 of inst : label is "5A5964949D924B72342E4B108208D64FA592A3750B92C4A0823593AB90CE4A41";
    attribute INIT_11 of inst : label is "57CE8195C3A46523665CA6D6B853D2E2BDE2B958A23929075F49E7236775D511";
    attribute INIT_12 of inst : label is "6E552F94261575A6144F944995FD099099E59796695D9C8DF54D365237557C52";
    attribute INIT_13 of inst : label is "33A9F2738185D04B44840151939997976909A58A9464E665E550995193999794";
    attribute INIT_14 of inst : label is "80C8EB96979A574B86895909D464E7A42555D2A8A295B4BDE3207BA28A543B36";
    attribute INIT_15 of inst : label is "A73B82FF9A6D000000007585D92E6137A235E6D9B4BF74E39C953A62DCE251D0";
    attribute INIT_16 of inst : label is "D6106763634235B71955424E4A424E674324E6763C68D8D88DDDC2E6B47E79AE";
    attribute INIT_17 of inst : label is "9761CAE710939290758727618DEA35B7197195E69C739B81C8D5534BF94E4A41";
    attribute INIT_18 of inst : label is "0000000000001D4D77A2DDA36DC65C6579A71CE6E0511634089C236084235926";
    attribute INIT_19 of inst : label is "5753619999B7DA373C224D2612B3BB9B4BD99F6E766B87924A5B753F96DB4000";
    attribute INIT_1A of inst : label is "3511676494526261C15B716F08084455927F4A8941066675656D45517756B841";
    attribute INIT_1B of inst : label is "459D9269741CF158518AE6F74B868DB991115649855961462B9C6236B2978575";
    attribute INIT_1C of inst : label is "2211262EA61075F79D824727709CF3195E69C6549E79A54BFFE55D2E1A36E644";
    attribute INIT_1D of inst : label is "E6B56537528227E692D3A9C2E080B5266167D2A75266154A086966EF8A942833";
    attribute INIT_1E of inst : label is "98DC26369D65766D2257F5FD394198D296D693527D79CB98211C59CB9CCA427A";
    attribute INIT_1F of inst : label is "A72349CBCA234992584B77741CA2379973713489CB265054C87BF1C232E59C24";
    attribute INIT_20 of inst : label is "54DC72C9941533288D66722798489201CB9142E9C8D249B72361C650418A12B9";
    attribute INIT_21 of inst : label is "426146A7292610D7F465A49E5B185E5637D2497263526DC8D84932C9612DDDD0";
    attribute INIT_22 of inst : label is "35E4AD92561EACF5985CF081F48DCF089453B82759715FF5D65945163D2E7676";
    attribute INIT_23 of inst : label is "51E690298092E49B4A4D09F79C6274B234A615819B4A099A4D282649F59E6352";
    attribute INIT_24 of inst : label is "000000000000000000000450CAAAAAAAA000000000000000000000022213FC65";
    attribute INIT_25 of inst : label is "499F4B5264A46427528557243081104104104104104104104104120820800000";
    attribute INIT_26 of inst : label is "674133EF9A52B6E15139B8944666257D85554D28227D2E4A4392C49934A02E7D";
    attribute INIT_27 of inst : label is "9C2E713D24E4A4645893A53FA525A73053A73CF7E79FED9B7988D66BFBEB4545";
    attribute INIT_28 of inst : label is "1C152347163260D934BF4394E91430730CF949E47A919B6423635F6242342413";
    attribute INIT_29 of inst : label is "725A6D908550227A590750227279863478D69B64657F7DF7DFDD65190F7A6624";
    attribute INIT_2A of inst : label is "5279C6485551A594CA46424E5D282079CB5266D282039CB52661B67927D891E2";
    attribute INIT_2B of inst : label is "291919E7B92E6A3723728D7F3CF7E655728D6C71CF7D092929B66D64DA52901D";
    attribute INIT_2C of inst : label is "D94B2B6E9D37195E69E1567279A59CA35235652618561060897D892909390979";
    attribute INIT_2D of inst : label is "2192464B6CBD5090B9FBA9841071A2F080BB0B9CCE739D4990EA63499D8C1A8A";
    attribute INIT_2E of inst : label is "0750709792D5929B6DF5DB8AE22749982E638D3902086279AE7B192864BE0BF4";
    attribute INIT_2F of inst : label is "7B54450708674192D64939BB7B85CF081C493D67D84A624A427D2E676157DA59";
    attribute INIT_30 of inst : label is "1141C21BD40608677199246E173C2063C4B44AD19DCD73544507086F43D19DED";
    attribute INIT_31 of inst : label is "82612B3812397F4E0ECCE772E3975CACE5D72C3975CB9C997195E69BBE2A5285";
    attribute INIT_32 of inst : label is "679A5C6195D2655D92373C2279295126710E373C225924152C87FBFFE19E4A2F";
    attribute INIT_33 of inst : label is "8B30062CC3194C2E5B9AC65A499969657924E79E84ACEEE6D2F46B5D23AC32BB";
    attribute INIT_34 of inst : label is "EE6D4BD1A2DF26C5CA9575A5171A5D6DDA9672AA5553787EA5DE7FFC6C900001";
    attribute INIT_35 of inst : label is "F6373C22603000024098EEE4FDFFFFC654545433A3FBB5EA4CC8845CBDF15DDD";
    attribute INIT_36 of inst : label is "CBAB2058EEE51FEDE7794B1831CC9320931FA64F9B9892CB2D3EBFAF624F5FFF";
    attribute INIT_37 of inst : label is "1C0AE3A173C2261EFBE0E9162E6770F2675A61D577942CF1A65373FA49BF16EA";
    attribute INIT_38 of inst : label is "F49F4B689C59375764124945D554158EE43A5DF8F49CE75B174B976412A40C39";
    attribute INIT_39 of inst : label is "2575589549041BDC6E638969095055555E984356AE1AC5DDDD555149D05F6891";
    attribute INIT_3A of inst : label is "5463895941577D77D75A2F49BA99955E4E39E9225373C2079E84ACE26D9B8465";
    attribute INIT_3B of inst : label is "D9B8615E7E5D5705CF0896DA6D9B8518ACB04E5C9552C8FC9695044444561527";
    attribute INIT_3C of inst : label is "E5ADE65E59E4B54758754755517B29F5397A1A83685CF0894E4A4D4B855B5156";
    attribute INIT_3D of inst : label is "E62F71E58D5D61D51D55479C797273C236D39842CA079697DA073C236D39E4A1";
    attribute INIT_3E of inst : label is "EEC7B1170050B3B82D623822C0C999B305CF3CEF89CF8E3E8923787330FBEA44";
    attribute INIT_3F of inst : label is "1619094555737F368A0CEC9D55D58DCF081B5A33332488884DDDDC515150CF8F";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "758CB312B371CB0C30F1C5C5C1D1D00078DC33331020BA68A01C5D91C30E9D75";
    attribute INIT_01 of inst : label is "EAE0B382CEC1901C31FD7A5FAC93C7A1F5C0DFAFCF1DB999802E002187DD633F";
    attribute INIT_02 of inst : label is "8CFCFCCCECB5CF2C75C557CC8733332DCB5CF397C637D3C738F3CCC76EAE0806";
    attribute INIT_03 of inst : label is "874FC901901F72BA0ED51038480DD703A00C72E6131D7801223E33BEF0F79312";
    attribute INIT_04 of inst : label is "D52164C8783B5408CEEA1E041A405FA724064F101822221C7C901900F72B9958";
    attribute INIT_05 of inst : label is "2EA54350D4350C2820242C2190590490490490680398B00B00B00B00B020342D";
    attribute INIT_06 of inst : label is "242B51802E0809F41F775AAAAAC45F0645C43D30B8231B32E0BBFF7527D2283C";
    attribute INIT_07 of inst : label is "931E4A01E33C703913C02E08057901D1F013F428CDC1C1C8DE48A1FFE2DCFDDD";
    attribute INIT_08 of inst : label is "738FEDCEC1E7E507CA9FF5445DC3E70424C6711327AB253187E87EEE1A02879E";
    attribute INIT_09 of inst : label is "5CA30C00420831932D8B0D8B1E0737727CBD75CF5DF0B63B612E9E9C9C5C5C5D";
    attribute INIT_0A of inst : label is "8DE7204101804F77DCFF3FCFF3FFF70300007075C7C48C77175D7E7CC8126071";
    attribute INIT_0B of inst : label is "DBA61C73D77C17078764F0793709D2E89D2E92E9F278D1DB2C0D1DB2CCD1DB2C";
    attribute INIT_0C of inst : label is "44242849C04140A0F8F805108EF5937173707CBBC406E1A074E021D93C1D72DC";
    attribute INIT_0D of inst : label is "AB7D75D7B05DF6726707A7E737D2C9CC9CC9C85085485885C400020283CF0F01";
    attribute INIT_0E of inst : label is "94CB7D033CBADF92F8975E5DFB30A5F9C1D679D185D2C7D1B3CB4B076B6B7E4B";
    attribute INIT_0F of inst : label is "1F35CFEDB5B5D75D7873D77F8F5DF0BCCBB9F1CD4B532DF5073D0CB5EE7C7392";
    attribute INIT_10 of inst : label is "E1CF5DFE3D77C2F32EC7E7F02D4CB7E41CF832D7B1F9FE4A532DF80CFB05C5D7";
    attribute INIT_11 of inst : label is "E827A9FA09E47F32C6911FA4E00B8AD2C372C7A04217175C7CD73F36D6D75D75";
    attribute INIT_12 of inst : label is "F1A41DDC1C8DE71089C1F9C1F9001E71EF7D7B7B07927ECB23B2C9EB2C8E40C9";
    attribute INIT_13 of inst : label is "08F3F9B8C082B82E228A9E3A71717071F60703E3DC9C5C5C1C30713271717070";
    attribute INIT_14 of inst : label is "F3BF6F90FB7739E746B727274E5C1D1C1CD7E17237DEE048CF523848D7746E68";
    attribute INIT_15 of inst : label is "1D3F42A3B84C3221021093A27E13E89C4B2EBE7EA079F23EF69D9BDA3013F7B7";
    attribute INIT_16 of inst : label is "1FB016F2D2F12E9D7DF38DC5C5C5C1D6FB5C1D6FB86CBCB4CB99BC22E2390FB1";
    attribute INIT_17 of inst : label is "30C003BF03717175C7C016C04BB12E9D7DD75E5DFC01F1808CBCEDE55DC5C5D7";
    attribute INIT_18 of inst : label is "840C840C40C424F49FC98839E35F75D7977F027C60175F2D2F3FB2CAFB32D77C";
    attribute INIT_19 of inst : label is "793C078727BD4720B822277370302C6D075CC5C65C6E037781E9D7D3BA74C84C";
    attribute INIT_1A of inst : label is "C175CF5DF009EDC78DE9D7F0ADAF5D7977ECC262C087C6AFD8D7237132FDE010";
    attribute INIT_1B of inst : label is "D73D77C30C02B31EC0C3BF49F746CBDAFD75E5DF1C72FB010EFC332EC07E3793";
    attribute INIT_1C of inst : label is "000008CC04A5C7CE5BEFDE96EBF8ED75E5DF5D7973D77E875577A79D1B2F4BF5";
    attribute INIT_1D of inst : label is "7D737EDE7709CF5DF354874BF081F357D3DD79DF357F7DE42FB7FD300330A680";
    attribute INIT_1E of inst : label is "FCB6FF2FF4C09F881BE4010047AB74B87B73FDCFD71FC5FAB0AFDFE5FF2DEDFE";
    attribute INIT_1F of inst : label is "BE12E7D664B2D5FBE2071B22364B2C5F49901C4FC6BC48DA62F0C749B17D741F";
    attribute INIT_20 of inst : label is "D66C31AF12349992CB57F11DF2E47880C577C97F0CBFEF009EC09E7DC067E0A7";
    attribute INIT_21 of inst : label is "D9C78BFCBFFC7C5F8BC87D7DFEF1D5CD0C77D5C9D2EBC027B02775AF881C6C88";
    attribute INIT_22 of inst : label is "2EDE5801328436E18482E0881C482E088BD3F42930187E175F7DF7DE9797F1C9";
    attribute INIT_23 of inst : label is "B05DF2474B797E6DCFF73F5D75C12DF92C1E07EC7DEC8F7FF7B23DFF5F77D2C1";
    attribute INIT_24 of inst : label is "003081003081003081000C710AAAAAAAA00C8CC40CCC8404040C8843003385D7";
    attribute INIT_25 of inst : label is "D5F5E7357CDC5C1EF9037B1A4840CF2C70CF2C70CF2C70CF2C70C03081003081";
    attribute INIT_26 of inst : label is "4774651C03E50380B71718E5C5C618FB0378F7B09FD797EDE1F9FD5FDEC097DC";
    attribute INIT_27 of inst : label is "76BFF7401CDC9D12B2743740DC9C9C48D1BCC108FD321801CFECB47757475465";
    attribute INIT_28 of inst : label is "729D1AD49D9BEA7E6075C9F65FADC8CC710DE34D40747600B2F2EEC9D92C9C73";
    attribute INIT_29 of inst : label is "C9C1D806DF7ABCFDFFDE7EBCFDEF032D4CB0760141C042403E24C027662A9C9E";
    attribute INIT_2A of inst : label is "EDEF0BFDF780DFF52DCDEDC9E7B0B61FE7357C7B0B61F67357C7603F3BB27509";
    attribute INIT_2B of inst : label is "0707C7DCFF3DFD2E12CCCB00C108FFB3CCCB108008BB2727076037BF73E8FF79";
    attribute INIT_2C of inst : label is "B1C432D45B8D75E5DF871CF5CF1CF332E92C5C9C781F7DD0FFBB27B7B7971747";
    attribute INIT_2D of inst : label is "89F987D4A2E318D2DF6BCFCF3A4A5BEA52F62DF311D9FCD5F4B3D8275B623124";
    attribute INIT_2E of inst : label is "5C72084B773EF07BEF1EB62DA77AFD74B7D8CB478BE1C9F7FDEF9F147C462E22";
    attribute INIT_2F of inst : label is "AEC5D7802F8AE0D0B5DF9955F7C02E080E29B86BB1C1C9CDCDD797D6C71F31CF";
    attribute INIT_30 of inst : label is "75E02BE2BE802F8AF0D77E5F00B82034ECE200883DABAEC5D780AF8AE4803DAB";
    attribute INIT_31 of inst : label is "D0370300050A40001B983AF9A8CAD66632B7998CADD5F55F975E5DF4C00CCA69";
    attribute INIT_32 of inst : label is "F3794BEFBE4901B00120B822375BEC902F8720B8222E180A1E5EF7BB81ADEC19";
    attribute INIT_33 of inst : label is "3DA560F6998247EDC777BEF8240BE05137DC737FDC0C093A01DCABD41B5682F5";
    attribute INIT_34 of inst : label is "B1A04772AAF113024EB218AC858AC46F4EB1113AC49337C6AECD7BB86C755558";
    attribute INIT_35 of inst : label is "E720B82225555554955BBC720100000A38C80506164B403800000024C61A2AAA";
    attribute INIT_36 of inst : label is "8E6E301BBC79011D22A8472E9A8159A84A3131A76C0EC5145A9D69717124CEEE";
    attribute INIT_37 of inst : label is "019F28F00B82213D34D805257C6A23193A01F35083FEEBE43DA08C783432B39B";
    attribute INIT_38 of inst : label is "EC7CCD547FCF1F31FBC1CF420DEC8700D0BFA8D7CC546814E8076A3B417E319D";
    attribute INIT_39 of inst : label is "9F033C5EC45DBC34F1FBEF5717B10DDDE07CE07EB8054050FA8CF2C43D31E47C";
    attribute INIT_3A of inst : label is "3F1BEF56C475F79C7DFC92EF8079733ED8BCDE17D00B82337FDC0C00180E029D";
    attribute INIT_3B of inst : label is "80E03F36F6CCDF402E088E01D80E001C22E00A3D7B71E455FE172321038E0B11";
    attribute INIT_3C of inst : label is "CCCCCC8CC4CCFC23F03F03F900870A1CBDF48C695C02E088B1C1C1EE0235C8DD";
    attribute INIT_3D of inst : label is "EF12F7DC61EFC0FC0FE403BDD4300B8223B07DC4C00373CD4720B8213B07CCC4";
    attribute INIT_3E of inst : label is "2910F4F84017D26B6B36507027639FA1320065A186001B60C6B337C699986AEA";
    attribute INIT_3F of inst : label is "034707A378D0C0612545A4FD3711402E08CACE5555495555211110A321141859";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "C0520828C45A20A20A37434343735812B60F4BBB366D84216A1400C3CF3C34D3";
    attribute INIT_01 of inst : label is "0644CA2310483B86834CD28D1CA36853636CCD33CDA0580912284A3B0D301480";
    attribute INIT_02 of inst : label is "D24106810603609010400369E0A04192E0360A236C3368DDA1D368DD20244E46";
    attribute INIT_03 of inst : label is "450DD404A48D81C34700AB849DAF006A359E0A2C0C93866188149B730E0C0828";
    attribute INIT_04 of inst : label is "003426529D1C02E60CF7808090128D2F50128D5891358D164D404A78D81C10D3";
    attribute INIT_05 of inst : label is "586BC7F1FC7F1D61616D6968510510510510510D6702856856856856856A9D15";
    attribute INIT_06 of inst : label is "10B089EE288EE34AF993E2CCCC46EF8CC563BFA8A23AA0C2CAC8304333F9856A";
    attribute INIT_07 of inst : label is "60A0AB035334D9E360EE288EE4562174F9A8CAB24343436A64ECF933CF433E09";
    attribute INIT_08 of inst : label is "D3133C33C34DD985E75CDA9A962355400D64BA0033F4310BCBC45CCC9D468AE9";
    attribute INIT_09 of inst : label is "0E7BE78EB8EB338A0693D293C00D0DA0D33CD35A249968088204343434343434";
    attribute INIT_0A of inst : label is "A654A6638A2A900301CC730CC330D09E9820D0D74740CC301D75DC77AD019850";
    attribute INIT_0B of inst : label is "EC2034A35D769D0D1D29D1D04B8360443604A04358D2434B066434B06E434B06";
    attribute INIT_0C of inst : label is "E64EF2CEC8687BC9A5A44B9925088991D0D0D8191E2B0A01D2C8874A74768100";
    attribute INIT_0D of inst : label is "7336034D712490D90D0D3340C340434CC0CC0004444884CC444000EF269A5A12";
    attribute INIT_0E of inst : label is "0241368335F4CD07340D3524990983766149DCE9C3704DE9D441010DFF33347F";
    attribute INIT_0F of inst : label is "7506592D11134D34D55549245A2499624184D430450904D81556441361350C11";
    attribute INIT_10 of inst : label is "5555249168926589069344C014241368555B104DA4D130440904D80CDA07475D";
    attribute INIT_11 of inst : label is "6033CCD81CF7349063B0342C089A2B4CF44CF083A31D1D75D41964B4444D34D3";
    attribute INIT_12 of inst : label is "486614C036A65496A094D094D2AA5E45E01C70030DB2C2C3BBA24B0B0EAECE03";
    attribute INIT_13 of inst : label is "49F680C9C9230A4CAA17BC95DCD0D0D3530DA973C274343434D0D895D4D0D0D3";
    attribute INIT_14 of inst : label is "EA6229B8D0039773A70D0D0D363434343669111331C1A862FDB7BC0CC30E4443";
    attribute INIT_15 of inst : label is "348CAB808000221119990498DD116A34090434DDA853633CD534A3664223626A";
    attribute INIT_16 of inst : label is "76408450506904828A2427474747674447767444B274181E818A99248A998DA0";
    attribute INIT_17 of inst : label is "D74123371DD1D1D75DC8844281A204828A0D35249C4CD8C1641907600C07475D";
    attribute INIT_18 of inst : label is "000CCCC48848812A34C82A3364A2834D49271336304D3504FF68505FF4904925";
    attribute INIT_19 of inst : label is "D04B8D0D0DE383A8A23A8DF909E9A65B852EE363363C88030348209082080CC0";
    attribute INIT_1A of inst : label is "88D35A249043434D23482890FCCF34D49264261B023363104264A993B904C8B8";
    attribute INIT_1B of inst : label is "4D68925D741188290223364741A74195DCD3514575DB24288CDEB90680DA0D04";
    attribute INIT_1C of inst : label is "04042E6EA2875D42113748445DD2CDD7565934D55549244500301DCE9D065773";
    attribute INIT_1D of inst : label is "340C3434D331DA2491740D233AD8CC034D04D004C134D348CF49259A23CA8BC4";
    attribute INIT_1E of inst : label is "D4133504D136377E114AAAAA0D1DD410D0D4D3534D4D04DB34B30D00D8034361";
    attribute INIT_1F of inst : label is "55A04C43449040D20D800D700449040D2AE4751D57236006BC284231D5345074";
    attribute INIT_20 of inst : label is "06B915C8C801AD0241135554DC055D405412310D241348D8847675D74233D995";
    attribute INIT_21 of inst : label is "534D7334CD34DA76403255500F03476765D34253604236211D8C50C8360035C0";
    attribute INIT_22 of inst : label is "043322A3986732C9CEA288EA80EA288EAF18CAB04D88D90D34D34D354D134343";
    attribute INIT_23 of inst : label is "7124950D3C513403434D0D34108844D504349D91D34CFD134D33F44D35135079";
    attribute INIT_24 of inst : label is "0810410400000030C30C30C30000000000044C956EA222044000088B0032434D";
    attribute INIT_25 of inst : label is "00D350C1353434350889904D0D400410410000000C30C3082082080000002082";
    attribute INIT_26 of inst : label is "FEECEDD7E3438A2202458C009163026489924D33134D13435CD1300D34CD1343";
    attribute INIT_27 of inst : label is "D3375DD0B47437BB80DD1DD0743437CE1A374F3C83CE22A34D281ECFFFFFDDFF";
    attribute INIT_28 of inst : label is "D134807074A754DDD85B5AD6ADE30E34C30B30F300D0D8A980604903488436D1";
    attribute INIT_29 of inst : label is "434362A534D33DA24934D73DA24906070010D8AB034000040001360D20AC3474";
    attribute INIT_2A of inst : label is "524977734D49249E034343435D33334D00C135D33334D00C034D8A8C7240DC07";
    attribute INIT_2B of inst : label is "2D2D0D01CC700C07807481E34F3C828F3481E38E38240D0D0D8A8D74D75DDCD3";
    attribute INIT_2C of inst : label is "1741B87421C0D35249ADB5A965A69D205404B434DA34D34DCD240D0D0DCD2D2D";
    attribute INIT_2D of inst : label is "4CD8335676C88EDECDF0CD34DD0F17040EC1DCDD034CD304D633740D21D0D025";
    attribute INIT_2E of inst : label is "B6D08420079240DE34838E6F9BBC045F7374810D37134340300DCD8B356BEC99";
    attribute INIT_2F of inst : label is "45A34DC8FF71A8D96249F08B4AD2288D219CB27243474353534D03486DB50A69";
    attribute INIT_30 of inst : label is "D3723FDC61C9FF7188C9242B48A234A0008AA68E6A1645A34DC8FF71BC8E6A16";
    attribute INIT_31 of inst : label is "FB909E9A2BB8AAAE11107C10C9DC147677051E9DC140D40D0D352496688F20B0";
    attribute INIT_32 of inst : label is "F8C0AC38D3D05AC1E3A8A23A8CCD3907B0ABA8A23A8C051A2B8B1B3309C00C80";
    attribute INIT_33 of inst : label is "D54A8755251CEA730007C34C416D31078CCEB803427A6997614E7E2CEC11CCC8";
    attribute INIT_34 of inst : label is "08368039D78B1958C707B4C1E34C1E38E707B15C1E361BDDC086333272BAAAA1";
    attribute INIT_35 of inst : label is "CBA8A23A800000002A114550000000038A14576434D41A0C5010100C6DB4B333";
    attribute INIT_36 of inst : label is "2F0C789145535B155A7A854DACDACACB834B5120812CEBAEB8752B5B51692CCC";
    attribute INIT_37 of inst : label is "0ACFACFA8A2398DFBEFD90F0723AB7B03A837840BACDEE7A3614046C22034BC2";
    attribute INIT_38 of inst : label is "40050514730D3CC377614702EED41995F3BF2A0B50069B434B83DA97A11748AC";
    attribute INIT_39 of inst : label is "374B963D413DCF433C0BCD0F0F506E66C0DE08DE322000E49326F541B0D3403C";
    attribute INIT_3A of inst : label is "4C8BCD01419B5D75D34C904F80D0DB9F38BEFD11EA8A239803427A60A2AC8834";
    attribute INIT_3B of inst : label is "2AC8B090202666EA288E6E0362AC89CEB288A79CD5914000DE0D333332264504";
    attribute INIT_3C of inst : label is "C0D2C12C1AC0FD4B44B46B48520A4C35CC008D0A4EA288E63343434C88992A66";
    attribute INIT_3D of inst : label is "F2907C30034E12E1AE214BCF102A8A239B8CD427A64803538398A239B8CDC0D6";
    attribute INIT_3E of inst : label is "5078355480095010858896926955151504D94D1760D95345E0261BD431351C09";
    attribute INIT_3F of inst : label is "234DCDB992665A4313291CDF995829288E5160000002222200000028515D90D3";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "701C32E40B00C33CF1F0C0C0C0E0F43002C20333F034D0181806A671C71C1C71";
    attribute INIT_01 of inst : label is "707801D02C01C400F1C030870021CF01E0C0C703073D01C1E0078101C31C070C";
    attribute INIT_02 of inst : label is "0072C072C030C32CB2E101C7871CB02C030C31E1C731C0C71CB1C7C307078030";
    attribute INIT_03 of inst : label is "0187C1102E07000F30F033000C0100D2F0047FF40D1FF0C0331FFF1CBC0702E4";
    attribute INIT_04 of inst : label is "C30018F0FCC3C082C31E1FC01C20C7C3044087C01E0C34047C1102C07000EC3D";
    attribute INIT_05 of inst : label is "5CCC0C03C0E0371FDF9B5B1803003C038034033C010CBC0BF0BE0BD0BC18FCC2";
    attribute INIT_06 of inst : label is "081CD41007410F4FF4CDF03333434103C13034401D043CF0750F0C3003453379";
    attribute INIT_07 of inst : label is "031F9CC0F31C352FC35007410C10404CD500CD4FC0C0E0DCFF74230F0230F35E";
    attribute INIT_08 of inst : label is "78E0F10F00C7420114CC73321C41C0003D340300037003073370133350C001F0";
    attribute INIT_09 of inst : label is "61461861451008733CB31CB31F03031C303471DE1C7573C73F3C0C0C0C0C0C0C";
    attribute INIT_0A of inst : label is "8FCB61C043DC1CB02C0B02C0B02C0F4240003031E1C00C07031C731EDC00201A";
    attribute INIT_0B of inst : label is "07071CC1C71C0303C3087C3CF200F3C00E3C13C0C03FC0C13DCC0C13D8C0C13D";
    attribute INIT_0C of inst : label is "CF3C906F40F032407070073CFCB073F0303038F1C101C1F0307430C21F0C702C";
    attribute INIT_0D of inst : label is "C31C71C7301C7030030302CC31F3C0C4400404804804804808C003C901C70701";
    attribute INIT_0E of inst : label is "304F1CB31FFCC7A99AC71C1C7C7531D0404C7B3400F3C734038F8F030F031FCF";
    attribute INIT_0F of inst : label is "1C71C704FCF0C31C7071C71C1E1C75704F0CB30CC0C13C73C71CF4F0C32CC330";
    attribute INIT_10 of inst : label is "C1C71C707871D5C13CB2CC300304F1C71C71D3C32CB30CC0C13C71CC72C0C0C7";
    attribute INIT_11 of inst : label is "C30340B0C0D02C13D00C0FC37401DC50C750C70CD003031C71C71C13E3C30C71";
    attribute INIT_12 of inst : label is "D10C061F0D0FCB710DF87DF87F03CC7CC71C7CB0030C304F530C30C13D4C31C0";
    attribute INIT_13 of inst : label is "01D79341C0103137701123FC34303031CDC353031F0E0C0C0C7C353C38303031";
    attribute INIT_14 of inst : label is "C8888F107CB0F1ECD00303031C0C0C0E0FFFC000301C100DC10E7000C07CB7FF";
    attribute INIT_15 of inst : label is "0C0CD40C700022222222CF307401CC1CC13F1C743011E030700C21C0B431C840";
    attribute INIT_16 of inst : label is "1C3333E3F3C13F2C70CBC0C0C0C0F0F3C30C0E3C1D08FCF04F3101CF7730071C";
    attribute INIT_17 of inst : label is "71C8031F84303031C7C013C0CF3D3F2C70C71C1C7F00B40404F2F1CC01C0C0C7";
    attribute INIT_18 of inst : label is "CCC888888888B3C41C01DC01CB1C31C7071F802D02071E3C0D7833C2D013C71C";
    attribute INIT_19 of inst : label is "3CF10303033D0D401D04071CF424344101B5C1D01D0B40B0C0F2C32C7CB3CCCC";
    attribute INIT_1A of inst : label is "2071DE1C7000C0C300F2C70C3C0D1C7071F1D403C802D0CB0FC373FC70B0F430";
    attribute INIT_1B of inst : label is "C77871C71C00C7F0CC031C31CCD0CF0CB471C1C71C73C3000C7F013CF031C3CF";
    attribute INIT_1C of inst : label is "040419955531C71FCF02DC23C0B07471C1C71C7071C71F010007C7B3423C32D1";
    attribute INIT_1D of inst : label is "2CC31F1C70035E1C704F03043501C331C71C732C331C71C00D071D1003000D84";
    attribute INIT_1E of inst : label is "78F02F3C73C01D0001FC0F03030C38F03C7871E1C7877C70FC20C74C71C0C0C3";
    attribute INIT_1F of inst : label is "1C13C74D4C13CC72C201A59C74C13CC7C2731CC74D2C81F093CF6703531C740C";
    attribute INIT_20 of inst : label is "F09CD34B307C25304F31D32C73CCB4004CB7034704F1CB1013C41C70C0034507";
    attribute INIT_21 of inst : label is "C0C3031C0B1C3C0C70C81C72C0B0C0FF0C71C3C0F3F2C404F107134B08069671";
    attribute INIT_22 of inst : label is "3F1D2DC8701C0077010074100C10074100C0CD4CF00031C30C30C30C0731C0C0";
    attribute INIT_23 of inst : label is "301C700308B31D31E1C7871CB5C13C023C0C030031C03CB1C700F2C71CB1F3C1";
    attribute INIT_24 of inst : label is "0410410410410400000010410000000000000C000C00000000000003003071C7";
    attribute INIT_25 of inst : label is "CC71CC331C0D0E0CB043FD3C00C0082082082082041041041041082082081041";
    attribute INIT_26 of inst : label is "2223202C41F043D0C7CB4031F2D00FC743FFC70031C731C0C0B30CC71C0231D0";
    attribute INIT_27 of inst : label is "3031C30C0C0C0C70F030C30C0C0C0CF2C21CB3CB0CB1FDC1C704F10010103322";
    attribute INIT_28 of inst : label is "300C13CB0C21C0742011C0B0873C72CB1C73CB2CB0303F7013E3F1C0C13C0C30";
    attribute INIT_29 of inst : label is "C0C0EDC01C7035E1C71C7035E1C7023CB8F03B70B0C000000033C00307700C0C";
    attribute INIT_2A of inst : label is "C1C702D1C7081C72C0C0C0C0C70030874C331C70030874C331C3F70B0C7032C0";
    attribute INIT_2B of inst : label is "0303032C0B02C33C13CB4F3CB3CB0CB1CB4F0CF3CBC7030303B7071C71C0B471";
    attribute INIT_2C of inst : label is "F0C013CB4F1C71C1C7C71DE1C71C72D3F23C0C0C3C0C30C0C7C7030303830303";
    attribute INIT_2D of inst : label is "00B302CD807611D1C70CC71C7C02384001C02C72C0C0B0CC7031C303CF0C7004";
    attribute INIT_2E of inst : label is "1C70000CB02C7033CB0C32ECBBB0D07C71C3CF030700C0CB02C00B302CD80760";
    attribute INIT_2F of inst : label is "0DF1C7000D01C0F571C70CD1CC60074200701DCC70C0C0C0C0C731E3C71C71C7";
    attribute INIT_30 of inst : label is "71E00B4070000D01C0C71F31801D080B3F7714C37B370DF1C7802D01C3C37B37";
    attribute INIT_31 of inst : label is "040F42400043C0D0EDFF70D341F0F4D07C3D341F0F4C74C7C71C1C74400C0CDC";
    attribute INIT_32 of inst : label is "1C70F2C30CC0D33F00401D040780CC0C0B09401D0434030007DD4CCCE532C01C";
    attribute INIT_33 of inst : label is "40000D000037C901C0B02C300340C00E07089CB03D090D10806143F6F53040CD";
    attribute INIT_34 of inst : label is "D108C185007300D3C03E370F8F70F8C7C03E3040F8F18C440F638CCD47D00003";
    attribute INIT_35 of inst : label is "3D401D0415555555404000055555555C7C300F0B0F4030031010103C0D37CCCC";
    attribute INIT_36 of inst : label is "C0B70400000F33070F04C18027C00243D3034004C34470000035C343400B4333";
    attribute INIT_37 of inst : label is "000D00D401D0407C30CC0C20450730100700C3C0720222C81FD7DBEC104CB02D";
    attribute INIT_38 of inst : label is "1C10C1CCB0C71C31D0800701CFCC0FC0CF3D1C4D0C30870107030710801F0024";
    attribute INIT_39 of inst : label is "0C7FFC0CC00C0C7031C3C70303303FFFF030C031DD0000AA54FFE0C03071CCB7";
    attribute INIT_3A of inst : label is "F203C7C0C0F1C71C71C013C070303FF2C03FC401F401D040B03D09003DCB400C";
    attribute INIT_3B of inst : label is "DCF407F2F2DCFF10074101C0EDCF400D007410FC33F04E9871C3222222FF3300";
    attribute INIT_3C of inst : label is "0C300F00F80C00D03C03E03434CC831E51C00C0205007410C0C0F0F743F0DCFE";
    attribute INIT_3D of inst : label is "2F13C71C30F0F00F80D0D0B1F02401D040FC33D09000B01D0D401D040FC30C30";
    attribute INIT_3E of inst : label is "00C0080000000000000000000000000003C0B7C103C02DF043318C4B13D040CC";
    attribute INIT_3F of inst : label is "00030373FFF0C0B0000BC4723FD010074100015555544444555555F0C03C2C3D";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
