-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(12 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S2
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (1 downto 0);
      ADDR  : in  std_logic_vector (12 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (1 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(12 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(12 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_01 of inst : label is "FFFF0000FE7D4C4CAA55FE7EFFFF00003FFCEEE055AAAAFD2D5F0AA02F580AA8";
    attribute INIT_02 of inst : label is "F000FC000000000007FF55552DEF00A87E7D4C4C1FFF00002FEF005410001FFF";
    attribute INIT_03 of inst : label is "F000FC00FFFFFFFFF547FFFFF800F000FFFFFFFFF457FFFF00000000FFC0FFFF";
    attribute INIT_04 of inst : label is "FA0F000F000F000F002F000FC0FFFFFFF01510FFFFFFFFFF1FD1FFFFFFF0FFFF";
    attribute INIT_05 of inst : label is "0A8001F0001400F20000000000000000008000000000BF4000000000000F000F";
    attribute INIT_06 of inst : label is "0BE0000000001680F00FFFFFF000F003F000F014F000F0000F00FFFF3C3ECF80";
    attribute INIT_07 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF0003000301500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "5000FC00900000000000C000F410FFF00000555501F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "0000001E0000000000000000B02F0000001503FF03DF0000000001FBC0FF4FFF";
    attribute INIT_0D of inst : label is "800000000000C100000300000AAA00010FE703FFDF900000AA00FAC0FFD6FC00";
    attribute INIT_0E of inst : label is "00000000AA800000008300000AAA0001FF802000AE00FFC083FF0020000401FF";
    attribute INIT_0F of inst : label is "E0FF0FFF5500FF00000000000AAA000000000000AA800000000000000AAA0000";
    attribute INIT_10 of inst : label is "0004FFFFE00F000FC00F800F8000000F002FD00F000503F7B0350000000503F5";
    attribute INIT_11 of inst : label is "800F0003000F0000003F003F02FF000F00403FFFC3FF0000FFFFCEAA8BFFFFF0";
    attribute INIT_12 of inst : label is "FFF3C00FA50F9A0F042FBE0FFFFFFFFF000000000000000000000000C00F800F";
    attribute INIT_13 of inst : label is "0FAB0000005E002C0000003ED2AB0000FFFFFFFFAFFEAAAA0000ABEAFFCF000F";
    attribute INIT_14 of inst : label is "FEFFFFFF0FFF000000FF0003FA870000AFFA0000E80F0007FF0FC00F002B0000";
    attribute INIT_15 of inst : label is "FFFF8E385D75FFFFFFEAFFC4BBFF23FFEB7FFFFFE7CFFF7FF3B3FFFFFF57FF57";
    attribute INIT_16 of inst : label is "E0FF57FFFF0BFFD5D803FFFFFEFFC97FFE29FF5F68BFF5FFFFBFFD63C027FFFF";
    attribute INIT_17 of inst : label is "0000005F000300005D60FFC4FFEA8E04197523FFBBFF8238FCBFFFFFF93FFFFF";
    attribute INIT_18 of inst : label is "056A002AA950A80000170FFFD400FFF000FF0002FF0080000000F500C0000000";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4FFFC0007003FFFE080004EFF0282";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFF5555FFFF00000003";
    attribute INIT_1B of inst : label is "0009C009C0090009600060036003600000005500000000550000666600006666";
    attribute INIT_1C of inst : label is "0003000300030003FFC3FFC300030003C000C000C000C000C3FFC3FFC000C000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000555500005555FFFF55550000555500005555";
    attribute INIT_1E of inst : label is "0000000000004000000000010000400000000000000000010000000000000000";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFF2FFFFFFFFFF800000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0033000F0000000AC04395BC0000D5E800000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "00CD00CC00000000735C330C00000000005700C00000000035C030C000000000";
    attribute INIT_23 of inst : label is "00CD30CC00000000735C330C000000000D4D00CC00000000735C330C00000000";
    attribute INIT_24 of inst : label is "01D60000000000A000000A00974000000000029C004000003FD8000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "CD73CC03000000005CD70CC30000000035CD30CC00000000735C330C00000000";
    attribute INIT_27 of inst : label is "3703303300000000373733330000000017350303000000003737333300000000";
    attribute INIT_28 of inst : label is "000F000A00FF0000F000A000FF00000000000FF5000000000BF03FFC00000000";
    attribute INIT_29 of inst : label is "0055055500150000550055505400000000550555001500005500555054000000";
    attribute INIT_2A of inst : label is "30DC30CC00000000DCDCCCCC0000000003373333000000003737333300000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "00EF1F400000D000F8000FF80150000001AF1FF50000D001F8001FFE01500000";
    attribute INIT_2D of inst : label is "00000000000000000000000000000000C07CE000FFC9FFD53D03000B63FF57FF";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "008F003F003E00004C00FC00400040001310054B00000000AEA0FE4005000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000800000000";
    attribute INIT_32 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000003";
    attribute INIT_34 of inst : label is "000200FA00000000A800BC0000000000000A00FE00000000A8003C0000000000";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000009000000000000000000000000";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFCFFFCFFFC";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "003F02FF005F0000FC00FF80F500000002A20FFF00000000FFC0FFF41D000000";
    attribute INIT_39 of inst : label is "E100FD22F804D7FD00BF206B042F7F57E0038000D34FD7FD08A71882E02B7FFF";
    attribute INIT_3A of inst : label is "0000000B000000002800FFE01F4000000000000000000000000002003F500000";
    attribute INIT_3B of inst : label is "03FF02FF07F4002AF800FFF00000800000FF03FF00050000F800FFF040000000";
    attribute INIT_3C of inst : label is "00FF0FFF00170028FF00FFF0D400000000FF2FFF00050000FF80FDD0FD000000";
    attribute INIT_3D of inst : label is "03FF3FFF017F002AFFC0FFFCFD40800003FF3FFF005F0000F3E0F7F4FF40A800";
    attribute INIT_3E of inst : label is "1FFF17FF11B40002FFF8FFFC000000000BFF17FF01B40002FFFCFFD000009A80";
    attribute INIT_3F of inst : label is "0EFF003F007F0282FFE0FFF0FF4022004EFF003F00070696FFE0FFFCFFF48000";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_01 of inst : label is "FFFFFFFFAF3CF9FEFFFF513FFFFFFFFFFF7C2AF8FFFFFFD01EAD001E1EA430AF";
    attribute INIT_02 of inst : label is "0000F400FFFF00000007FFFF3FFF0B57FF3CF9FE0FFFFFFF3EBF0B57FFFF3D15";
    attribute INIT_03 of inst : label is "0000F400C5F0F6FFF000FFFFFFFFF000FFFFFFFF0000FFFFFFFF0000FFC0FF80";
    attribute INIT_04 of inst : label is "EC0F800F000F000FFFFD000F901FF60BF000E0FFC3FFFFFF0000FFFFFFF0FF50";
    attribute INIT_05 of inst : label is "57C00000000000F5FFFF0000400000000BF0000000005400FFFF0000000F000F";
    attribute INIT_06 of inst : label is "BFF4000000000040F003F47FF00BF000F000C000F000F000CF004BD0C7EDF1E0";
    attribute INIT_07 of inst : label is "55555555D555D55555575557AAAB000300000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "0000FC00C000080003F01800F000FDA0000000002ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "000000010000000000000000C0FF00000000003B03C318A000000245C03F0FFF";
    attribute INIT_0D of inst : label is "C800000003F00000000300180FFF00020FD0017FC3C0A008F000071801E0FF00";
    attribute INIT_0E of inst : label is "00000000FC000000001B00000FFF00005AD8C000F00007001B4A00E000000007";
    attribute INIT_0F of inst : label is "F03F0FFF0000FF00000000000FFF000000000000FC000000000000000FFF0000";
    attribute INIT_10 of inst : label is "FFFBFFFFD00FC00F000FC00FF00B0005FFFF400F00000000C001000000000020";
    attribute INIT_11 of inst : label is "F00F000B000F0055000F003F0FD7002AFEBF07F7C1FF157FFFF0EFFFED7FAAA0";
    attribute INIT_12 of inst : label is "C013C0073C0FCF0FFFFF1C0FFFFFFFFF0000000000000000000000000003C00F";
    attribute INIT_13 of inst : label is "0003000300FC003CFFFF0074FFFFE000FFFFFFFF83C2C444FFFF555583CF028F";
    attribute INIT_14 of inst : label is "FFFFF27F0F020A8000030003BFFF000B03C00000FC0FFD53C00FC00F0035057F";
    attribute INIT_15 of inst : label is "FFFFAEBA1C71FFFFFFC4FFDD23FF57FFFEFFC9BFFEBFDAE7FBFBFF3FFFFFF57F";
    attribute INIT_16 of inst : label is "FAFF947FFFAFFD16C6BFFDFFFFFFE403FFEAFF07ABFFD0FFFFFFC01BFE93FF7F";
    attribute INIT_17 of inst : label is "0000000300AF00001C41FFDDFFC4AE98207157FF23FF06BAFFFFF63FFFFFFC7F";
    attribute INIT_18 of inst : label is "00002D4000000178000007F74000DFD003FF003FFFC0F8000000C000FA000000";
    attribute INIT_19 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5540FFFC0000000FFFF8FE0001FF56FB";
    attribute INIT_1A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFF4FFFFAAAAFFFF00000003";
    attribute INIT_1B of inst : label is "0009C009C009000960006003600360009999000099990000AA00000000AA0000";
    attribute INIT_1C of inst : label is "0003000300030003FFC3FFC300030003C000C000C000C000C3FFC3FFC000C000";
    attribute INIT_1D of inst : label is "AAAA0000AAAA0000AAAA00008000000000020000FFFFAAAA8000000000000000";
    attribute INIT_1E of inst : label is "0000000080000000000200000000000080000000000000000002000000000000";
    attribute INIT_1F of inst : label is "FFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000";
    attribute INIT_20 of inst : label is "003900000000002DE24B55400000B71E00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "00CC014500000000330C51540000000000AB00550000000030C0154000000000";
    attribute INIT_23 of inst : label is "2ACC104500000000330C5154000000000E8C054500000000330C515400000000";
    attribute INIT_24 of inst : label is "00150000000000F800002F005400000000003FE400000000016C000000000080";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "CEB34551000000000CC35455000000003ACC154500000000330C515400000000";
    attribute INIT_27 of inst : label is "3B1715110000000033331515000000002B3A1515000000003333151500000000";
    attribute INIT_28 of inst : label is "000300BF0005000FC000FE005000F0000FFA0000000000003FFC07F000000000";
    attribute INIT_29 of inst : label is "02AA02AA0000002AAA80A8000000A00000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "30CC105400000000CCCC5454000000002B331515000000003333151500000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "2FFD0000000005027F001FBD000080002FFF000000000500FF800BBC00008000";
    attribute INIT_2D of inst : label is "00000000000000000000000000000000C014FFD4FFFEFFE0140307FFBFFF0BFF";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0004007D0004002FBC0073C00000C0000FF4005500000000FD745A0000000000";
    attribute INIT_31 of inst : label is "0000000000040000000000001000000000000000000000000004000000000000";
    attribute INIT_32 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000003";
    attribute INIT_34 of inst : label is "003D0015000000005F00500000000000003C0015000000007F00500000000000";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000009000000000000000";
    attribute INIT_36 of inst : label is "FFFFFFFF5555FFFFFFFFFFFF5555FFFFFFFFFFFFFFFFFFFFFFFCFFFCFFFCFFFC";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "002F07FF0001002FF800FFD04000F8000FFF015100000000FFF8FFC000002E00";
    attribute INIT_39 of inst : label is "FFA0F004FEE8EA000A07440F2BBF042B4000C003EBBFC1701811100BFFFF9017";
    attribute INIT_3A of inst : label is "0000000000000000FE00FFF000000000000000000000000000000FE000000000";
    attribute INIT_3B of inst : label is "007F2FFF004003FFFF8055D00400F00002BF037F00000000FF80F4000000A000";
    attribute INIT_3C of inst : label is "03FF07F70000002FFFC0DFD00000E0000BFF11FF0000000AFEE0FF400000FE00";
    attribute INIT_3D of inst : label is "0FFF1FFB000100AFFFF0EFF44000FA002FFF13FF000000AFF7F8FFD05400FF80";
    attribute INIT_3E of inst : label is "1FFF2FFF000008BFFFFC5FD00000FA802FFF2FFF000000BFFFFC50000000DFF8";
    attribute INIT_3F of inst : label is "01FF00FF000502FBFFF8FFC05400FF4001FF000F0000A6FBFFF8FFFC5540FE00";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "007802803D540AA82AAD0AA81E3C002801F40AA8017E2AAA00F00AAA3C0F02A0";
    attribute INIT_01 of inst : label is "0000FFFFFFFFFFFF01FFFFFF0000FFFFFFFFFFF8FF40FFFF2D5F0AA02F580AA8";
    attribute INIT_02 of inst : label is "5F00FF400000700000000000BDEF03FF7FFFFFFF0000FFFFBFEF03FF74007FFF";
    attribute INIT_03 of inst : label is "5F00FF4003FF000002010A1500000017FF6F00005000DFCF140000A3FF340000";
    attribute INIT_04 of inst : label is "FA000000FE00A00000007F40300F00000600E068FFFD00000540577FBFC40000";
    attribute INIT_05 of inst : label is "1FDBFBF0D2BCFEF000552FFFAFFF0000FD1F03F82FFF000A4000E015FF800000";
    attribute INIT_06 of inst : label is "D00702F82FFF168A000F00000A80000307F40BFF03FF00BF0F0000003C3ECF80";
    attribute INIT_07 of inst : label is "FFFFFFFF3FFF3FFFFFFCFFFC0003000301500000006020002D5F0AA02F580AA8";
    attribute INIT_08 of inst : label is "3C1502AA3D5428000F540AAA3C0F2AA03C0002A83D5E2AA83C0F280A00000000";
    attribute INIT_09 of inst : label is "3C0F0AA83FDF280A3FFF280A0F000AAA3DE0282A000F0AA800F00AAA3D5F280A";
    attribute INIT_0A of inst : label is "3DDF280A3D1F00803C0F0AA800F000A02D540AA83C1F282A3C0F0AA23C0F2800";
    attribute INIT_0B of inst : label is "AAAD400FFE0080005AF0FF00000000000000FFFF01F82AAA0B5E00A00BF8280A";
    attribute INIT_0C of inst : label is "0000000000000000FFFFFFFC002FFFFE1EAA03FFFFFF0AFEE17F7FFFE000F000";
    attribute INIT_0D of inst : label is "FE0080005AF0FF00F0FFF00AF555FC7FF000F000FFFEFE8055FFFFFF000003FF";
    attribute INIT_0E of inst : label is "09000000557F0180F0FFF00AF555FC7FFFFEFE8055FFFFFFFFFF0AFEE17FBFFF";
    attribute INIT_0F of inst : label is "E100B000EAADF00FF000F000F555FC0030000000557F3000F006F000F555FC09";
    attribute INIT_10 of inst : label is "557FFFFFFE00A000F3C0FFC0E1FF03C04000FC001EAA03F50035FFFE1EAA03F5";
    attribute INIT_11 of inst : label is "E7D0003C003F02AA00FF00FF2FFF003F03D1FFFFFFFFAAAAFFFFFFFFFFFFFFFC";
    attribute INIT_12 of inst : label is "FFFCF550FFC07F801D00FFC0FFFFFFFF000000000000000000000000F0E0FFC0";
    attribute INIT_13 of inst : label is "3FFF005F03FF00BF00F002FFFFFFA800FFFFFFFFFFFF55550000FFFFFFF00000";
    attribute INIT_14 of inst : label is "FFFFFFFF3FFF000003FF555FFFFF002AFFFF5555FF00AAA8FFC0F50000FF2AAA";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFF83FFFFFF3B3FFFFFF57FF57";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "0000005F00030000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCBFFFFFF93FFFFF";
    attribute INIT_18 of inst : label is "0000000000000000016B3FFFE940FFFC03FF000BFFC0E0000000F500C0000000";
    attribute INIT_19 of inst : label is "FFFF0AFF3FFFFFFFFFFFFFA0FFFCFFFF0009DC77001800FFFFF8E800FFFF0BEB";
    attribute INIT_1A of inst : label is "F7AFFFFFDEBBF7FF0A1CD6278040000200000000FFFFFFFFFFFFFFFF00000003";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "003FFFFF003F003FFFFCFFFC003FFFFFFC00FFFFFC00FC003FFF3FFFFC00FFFF";
    attribute INIT_1D of inst : label is "FAAAF000AAAA0000AAAF000FF800FFFF002FFFFFFFFFAAAAF800FFFF0000FFFF";
    attribute INIT_1E of inst : label is "00000000F800FFFF002FFFFFF000FFFFF800F000000FFFFF002F000F00000000";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFF000F000000F000F0000FFFF";
    attribute INIT_20 of inst : label is "0033000F0000000AC04395BC0000D5E800000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "00CD00CC00000000735C330C00000000005700C00000000035C030C000000000";
    attribute INIT_23 of inst : label is "00CD30CC00000000735C330C000000000D4D00CC00000000735C330C00000000";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "CD73CC03000000005CD70CC30000000035CD30CC00000000735C330C00000000";
    attribute INIT_27 of inst : label is "3703303300000000373733330000000017350303000000003737333300000000";
    attribute INIT_28 of inst : label is "003000B507040FFA0E805E0010D008002FBC300AF0050000B60EC48307D50000";
    attribute INIT_29 of inst : label is "0155155501410154554055544140000001551555014101545540555441400000";
    attribute INIT_2A of inst : label is "30DC30CC00000000DCDCCCCC0000000003373333000000003737333300000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "000B05BF00000000E000F7E000000000000B055A0BFF0000E000E7E8D0000000";
    attribute INIT_2D of inst : label is "00000000000000000000000000000000C07CE000FFC0FFD53D03000B03FF57FF";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "003F00EF00FE00AAFF00FF80D140A5982AAB3FFF90000000F8F8FE901F400000";
    attribute INIT_31 of inst : label is "F63FF64FF3CFFF2AFC9FF19FF3CF3FFFFDA839FFFD9FFFFF445BFFFE9E5BFFFF";
    attribute INIT_32 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFCFFFCFFFC";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000003";
    attribute INIT_34 of inst : label is "0B9D3FF5007F00005BF07FF4F50000000BFE3EFF01760000FFF0FFE4F5000000";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE40AC0F6FE80FFFFA80FFC0B0AFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFF3FFF3FFF3";
    attribute INIT_37 of inst : label is "FFFF000000009999FFFF0000000099990000000000000000FFF6FFF63FF63FF6";
    attribute INIT_38 of inst : label is "007F03FF007F0000FE00FF80FFC0900002BF0FFF00010000FFF4FFF45D000000";
    attribute INIT_39 of inst : label is "E100FD22F83CD7FD00BF206B3C2F7F57E0038000D34FD7FD08A718A2E02B7FFF";
    attribute INIT_3A of inst : label is "000200BF00010000FF00FFFEFFF40000000000000000000000002FE0FFFD0000";
    attribute INIT_3B of inst : label is "0F2F2FFF7FFF0AFFFF90FFFE4040F82003FF07FF01FF0000FF80FFFAF480A000";
    attribute INIT_3C of inst : label is "03FF3FFF016B01FEFFC0FFFCE940800003FFBFFF005F0000F560F774FF40A800";
    attribute INIT_3D of inst : label is "FC00C000FE80FFD5003F000302BF7FFFFC00C000FFA0FFFF0C1F080B00BF57FF";
    attribute INIT_3E of inst : label is "7FFF7FFF77FD002BE406F8030540A0002FFFBFFF77FD002BA003F8240000E560";
    attribute INIT_3F of inst : label is "3FFF00FF01800BEBFFF8DDFC0090BB90FFFF00FF00180FFFFFF8DC770009E800";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "3EAF03C007A83C0F3EA8140F01FC2ABE0ABE140F1EAD1FA001F000F006B42D0E";
    attribute INIT_01 of inst : label is "00000000AFFFFFFFAAAAF7FF00000000FFFFFFFEAAAAFFF41EAD001E1EA430AF";
    attribute INIT_02 of inst : label is "2C00A9000000000000000000FFFF2F57FFFFFFFF0FE00000FEBF2F570000FF7F";
    attribute INIT_03 of inst : label is "2C00A90003FB00AA00700FC300000001FF3F00000000F1FA00008B75FFB4280F";
    attribute INIT_04 of inst : label is "EC000000FF00FF0000000000600709020070183FC7FCA80000000FC7FFC4000F";
    attribute INIT_05 of inst : label is "F7C57FE82FFFF4F0000007FF5FFF002A50032FFF857F02BF0000F400DFC0A000";
    attribute INIT_06 of inst : label is "00032D7F857F02FF0003007F074B0000000A3FFF005400BFCF004BD0C7EDF1E0";
    attribute INIT_07 of inst : label is "FFFFFFFF3FFF3FFFFFFCFFFCAAAB000300000000000606001EAD001E1EA430AF";
    attribute INIT_08 of inst : label is "07AA2D0F3EAA3C000FAA0F003EB43C1E07AD2D053EAD3C0F07B43EAF00000000";
    attribute INIT_09 of inst : label is "1EAD3C0F3D0F3CBF3D1F3C8F0F000F003C1E3EF4000F140F0AFA00F03C0F3C0F";
    attribute INIT_0A of inst : label is "3C0F3FBF3C0F0BF83C0F3C0F0AFA00F01EB4140F3EAD3EF41EAD3CBE3EAD3EA8";
    attribute INIT_0B of inst : label is "00000003FF00F800FC00FCF000000000000055552ABF1F800F0F00F03D1F1FBD";
    attribute INIT_0C of inst : label is "AAAA0000AAA80000FFFFFFFF00FFFFFF0000E02BFFFF3FFFFFFF1DBFFC00F000";
    attribute INIT_0D of inst : label is "FF00F800FC00FCF0F0FFF03FF000FF1FF000F000FFFFFFF80FFFBFE7000000FF";
    attribute INIT_0E of inst : label is "0000008003FF0013F0FFF03FF000FF1FFFFFFFF80FFFFFFFFFFF3FFFFFFF5FFF";
    attribute INIT_0F of inst : label is "FC00F0000000C003F01AF000F000FF0005800C0003FF4003F000F020F000FF10";
    attribute INIT_10 of inst : label is "0004FFFFFFC0F00043C0F7C0FC1403CA0000F0000000E0000001FFFF0000E000";
    attribute INIT_11 of inst : label is "FC000EB400BF03FF00FF00FFBFFF02BF01401FFFFFFFFFFFFFFFFFFFFFFFFFFA";
    attribute INIT_12 of inst : label is "F5FCFAA8FF403FC000007F40FFFFFFFF000000000000000000000000403CF5C0";
    attribute INIT_13 of inst : label is "155F2A8F03FF02FF000003FDFFFFFC0AFFFFFFFF5FF53BBB0000FFFFFFF0AFF0";
    attribute INIT_14 of inst : label is "FFFFFFFF3FFF3FFA015F02AFFFFFA83F5FF53BBBFF00FFFCF7C0FAA000FF3FFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFF51FFBFBFF3FFFFFF57F";
    attribute INIT_16 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_17 of inst : label is "0000000300AF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF63FFFFFFC7F";
    attribute INIT_18 of inst : label is "000000000000000000011FC30000C3F40FFF00AFFFF0FE000000C000FA000000";
    attribute INIT_19 of inst : label is "FFFF3FFF05FFFFFFFFFFFFFCFF50FFFFAA90400300010034FFFEFF8007FFFFFF";
    attribute INIT_1A of inst : label is "FFFBFB7FEBEBDCEFC12B81120202040000000000FFFFFFFF5555FFFF00000003";
    attribute INIT_1B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_1C of inst : label is "003F003FFFFF003FFFFCFFFCFFFF003FFC00FC00FFFFFC003FFF3FFFFFFFFC00";
    attribute INIT_1D of inst : label is "5555F00055550000FFFF000FFFFFF555FFFF555FFFFFFFFFFFFFF555FFFF5555";
    attribute INIT_1E of inst : label is "FFFF0000FFFFF400FFFF001FF000F400FFFFF000000F001FFFFF000F00000000";
    attribute INIT_1F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000F000F000000F000F00000000";
    attribute INIT_20 of inst : label is "003900000000002DE24B55400000B71E00000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "00CC014500000000330C51540000000000AB00550000000030C0154000000000";
    attribute INIT_23 of inst : label is "2ACC104500000000330C5154000000000E8C054500000000330C515400000000";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "CEB34551000000000CC35455000000003ACC154500000000330C515400000000";
    attribute INIT_27 of inst : label is "3B1715110000000033331515000000002B3A1515000000003333151500000000";
    attribute INIT_28 of inst : label is "03DC0B61037A00F0354049E0ADC05FC03005FF5E00000A28C843790500000BEA";
    attribute INIT_29 of inst : label is "2AAA0A82000000AAAAA882A00000AA0000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "30CC105400000000CCCC5454000000002B331515000000003333151500000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0AD60BFF000000009E8047B4000000000AFD00BF3FFD00007E00F7B000000000";
    attribute INIT_2D of inst : label is "00000000000000000000000000000000C014FFD4FFFEFFE0140307FFBFFF0BFF";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "00BF003D001D00BFFF007FF00000FE003FFFC7FF10000000FD7DFF0000000000";
    attribute INIT_31 of inst : label is "FF1FFD4FFEBDF7D6F4FFF17F7EBF87DF52FF1E54FFFFFE6FFFFD88A7FFFF6DA7";
    attribute INIT_32 of inst : label is "FFFFFFFF7555FFFFFFFFFFFF5555FFFFFFFFFFFFFFFFFFFFFFFCFFFCFFFCFFFC";
    attribute INIT_33 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000003";
    attribute INIT_34 of inst : label is "2FFE0F7A000000AFAFFCB9D00000FC8027FF0FFF000000AFFF7C7FD000006E80";
    attribute INIT_35 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03FF015FFFFFF506F03502FFFFF017F";
    attribute INIT_36 of inst : label is "FFFFFFFFAAAAFFFFFFFFFFFFAAAAFFFFFFFFFFFFFFFFFFFFFFF3FFF3FFF3FFF3";
    attribute INIT_37 of inst : label is "55FF00000000FFFFFF5500000000FFFF0000000000000000FFF6FFF63FF63FF6";
    attribute INIT_38 of inst : label is "02AF07FF000100FFFD00FFD04140F8006FFF0FD300000000FFF8FFD000002EA8";
    attribute INIT_39 of inst : label is "FFA0F004FEE8EA000A07440F2BBF042B4000C003EBBFC1701851105BFFFF9017";
    attribute INIT_3A of inst : label is "000B001700000000FFE0FFFD1F40283000000000000000000000BFFE7D400000";
    attribute INIT_3B of inst : label is "0FFFFFFF07F41F57FFF8FFFD2F00FCF80FF203FF00140BEBFFF8FFFC1050FC00";
    attribute INIT_3C of inst : label is "0FFF1FCB000100BFFFF0E3F44000FA002FFFF7FF000000AFFBB8FA905400FF80";
    attribute INIT_3D of inst : label is "F000E004FFFEFF50000F100BBFFF05FFD000EC00FFFFFF500807002FABFF007F";
    attribute INIT_3E of inst : label is "7FFFBFFF02506EFFE803F0240000F560BFFFBFFF037002FFE803F5400000F006";
    attribute INIT_3F of inst : label is "07FF0304001A8BFFFFFE4130A900FFD007FF00340001FFFFFFFE4003AA90FF80";
  begin
  inst : RAMB16_S2
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
