-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity cpurom is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of cpurom is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FB4D3B69A6C0C04A8D6098C1151AC1318A8D504DBA0850B2D405000000000109";
    attribute INIT_01 of inst : label is "8DFFB8E5CAA734412544B9358F8891B139B27B69E6DA46DE6F4D8FDEDB07E9F3";
    attribute INIT_02 of inst : label is "26375B8E4A862419EF8BFFE022B5A24AD461B8BAF2EEBB7A4F95386CE2A2C51D";
    attribute INIT_03 of inst : label is "42288884244A115457BD6919A449A4D98899DCD20999EB26E6C6641224D81012";
    attribute INIT_04 of inst : label is "039487D09840407DDE6EC635DA6C96AAD446B6EBFFD0A4440FAA9415EA020A02";
    attribute INIT_05 of inst : label is "D321A451BC829B6DBF67ED03E6189459B3D07A5F8F06101CC1338073128B95B6";
    attribute INIT_06 of inst : label is "599DEF3F56BB79E3A70A0F2C8490EDC395250EA93C545CAA2A25DF82545F6ED1";
    attribute INIT_07 of inst : label is "4E66723490EBFE329A93CDF70DF78E37843CFC586A367BCD70020001097B4433";
    attribute INIT_08 of inst : label is "FF2784291FC27F4E1C483DE9B6107A1A8EE5DC1F01E14D7CA9512A21009813E8";
    attribute INIT_09 of inst : label is "D0121E2A3F8FBEF8EEB371F373140F8B712E1F176090D00F1511FFDF7C7A4A30";
    attribute INIT_0A of inst : label is "511E33DF7DF631854C8F19191184A92A067FD0974008041383074961066C849E";
    attribute INIT_0B of inst : label is "7652D55556836C32C3663363C092E8814C98CB5A49A49EBEE895833FF99B6AF9";
    attribute INIT_0C of inst : label is "9533B2A44AA08229813FA49A492339E7E6E719D58AB90E63128D6E31B8D629A9";
    attribute INIT_0D of inst : label is "53A02162DD54B224729F6F546D5BDF12551F57A1FFC7C8F83CC486E10AA0822C";
    attribute INIT_0E of inst : label is "535115CD2AC84056B4DF3E99C37156F17E927E907EDB8E5C7524967989000000";
    attribute INIT_0F of inst : label is "A46D266766A0A92A0A922034035384AA11AEE5256A15C25AA319355954AB3735";
    attribute INIT_10 of inst : label is "27E1B4A01151FB3F07420283ED5212A42689548908E44000800200440000F44D";
    attribute INIT_11 of inst : label is "90D8654D144966555405268D2B9960A989D62A0C11520B90143F01C091260550";
    attribute INIT_12 of inst : label is "5A1FE35C51A7C7F1C58270438E8478C799A04A252D083DD936DF74B1CBE6755D";
    attribute INIT_13 of inst : label is "A440D5EE03D44A84381E6E5B039FBFFE4C2AF972E5157D42936DF8E1FFF55FF0";
    attribute INIT_14 of inst : label is "61308C56E091A3DC6371784555B6FCC1FF87AAC6FF4A7CBE2921FCCD965A1E01";
    attribute INIT_15 of inst : label is "3B649EDF19C8A2D0A4BB641BB64534E0059207D3B77D0FD885530D5AA3FD9C8A";
    attribute INIT_16 of inst : label is "8D760AA4A01785DF7339CC1D51B4393BFC8AE5476C837DEC8B4DA61FCD90ED93";
    attribute INIT_17 of inst : label is "022CA00115BB67FCA22DCC253C62E19C30842E4ADEDA6DD3E12E9334E1D5BAF0";
    attribute INIT_18 of inst : label is "1C692100E5E2B09FD7FC4A81412AB649D612CA7500CAF40038DCFE79CF1E7940";
    attribute INIT_19 of inst : label is "261987AD753861929030552500A997A5F8D5C5D5C521084CF202014A43744729";
    attribute INIT_1A of inst : label is "098455A06F2C910010912609C8846929EAE79FFDFFF8452528A8ACAC8A2A2A2A";
    attribute INIT_1B of inst : label is "A496466966D31D1E4198109A130779F981F61D0D098C86B990C93FDC4AFA1327";
    attribute INIT_1C of inst : label is "A67DB153168B55EBA366102D29BE3D950528A79DC7E9F0215088A55B3D868529";
    attribute INIT_1D of inst : label is "68930C97D94ECDBFD26583E330571012308479BFCD494B0A29112537CE348345";
    attribute INIT_1E of inst : label is "FCB0888219BE30D2E33F6B08B3493764E3D0E55B0E9EDC4980348D6147FA7E0C";
    attribute INIT_1F of inst : label is "D9453AB560C738000305510180075FAF8D54C2BC660046D5214D04A80C142819";
    attribute INIT_20 of inst : label is "00000800585810000010001010100048004800105D58351950709B1E10B25A42";
    attribute INIT_21 of inst : label is "AAAAAAA911000000000001104100000000000000000000000000100010000010";
    attribute INIT_22 of inst : label is "000000000000000000000556DF7FFFF80F802015031575030128000400040C02";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "00004000D304F2AB781E9DEB66EDC1B6AA25BE6D728DF1B2930E4D7BC5AC725E";
    attribute INIT_25 of inst : label is "9C47CB64C817B650E55AAD0D6DD2CD89770CE3A4DE023E6A954CCC28F9F80000";
    attribute INIT_26 of inst : label is "1B6D84AA70DB36C725EA954AA68496C9C464B7C96AA1BB0DDA5EA954AA684974";
    attribute INIT_27 of inst : label is "E9471A005561189CE0E5AA92809596C9E989996F020A954966849494B696AA42";
    attribute INIT_28 of inst : label is "6F6B7FB58524E45AE2ABFC37B8ADBFD4BFFBEB2D1BAA291BAD5968C37FA4DFFF";
    attribute INIT_29 of inst : label is "04AAE0844215DE8A2FFAAFFAAFFAB83D8E6F52F7E9825A09414B4DED2B550011";
    attribute INIT_2A of inst : label is "55C0A20618082A2288BC22AAA220AFBBAF7FECE0EAF796FECE4800000003E111";
    attribute INIT_2B of inst : label is "E1CF1A0EFFA2F66F62F0AEA08004155455551400100004000100C08202184405";
    attribute INIT_2C of inst : label is "000000000000000000F8A4FCEC262A12F1B77238D6C7D0F85302FF00000041F5";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "277C8B1F05550554550554155411677AFDFF0FF8FDFEF936FE9EF9AF23200112";
    attribute INIT_31 of inst : label is "D711353B01015151CDD051455054554044446622455514505010000040010541";
    attribute INIT_32 of inst : label is "7AB4980913011105141567313330333311EEFDFCFD6515545155515415500010";
    attribute INIT_33 of inst : label is "AD8D06B4037555555055551551DDC98100111015541572275554555511011550";
    attribute INIT_34 of inst : label is "00000000277775DDDDCFFF777731677BFDFFDFF8FFFEF9BFFFDFFDFFFFEFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "520366EE66939474AA7653B24034C0D30D30D30D30D3FFFF1D88BFFDE4E0DFF9";
    attribute INIT_39 of inst : label is "0BEF817D3F0FC0BF7E1C4E0458C0D2ABA02827E0936F6426DEC84A7653B2F9C1";
    attribute INIT_3A of inst : label is "F57F80632BA6813103B47B62A809B149E6A49C3524F2926949269000B49310B0";
    attribute INIT_3B of inst : label is "5BA5B0649567D669558937D2D4003042F03D7E80BBDBA0904FAA9D904948320B";
    attribute INIT_3C of inst : label is "DAD1AD68D6ADB35AD1AD6CD6B46B5B35AD1ED6CD6B7DFEF2F5AEB74B60965967";
    attribute INIT_3D of inst : label is "267249896ECC8080CC0F159F610A7ACB26D6366B5B3DAD1AD57B1B2F6B47B5B3";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000DBD9A747DB3C";
    attribute INIT_3F of inst : label is "2E00000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "8CB3068A215C2688400B33CA642092279AC8A24C88A28400FA01000000000181";
    attribute INIT_01 of inst : label is "13006A123459A75157236642634D1CC64067AFFEE9C85F412DA5C201E54232A3";
    attribute INIT_02 of inst : label is "11048728099D049B4A1DD513ECE8677C32C6155D74B557AA805A468008C9B920";
    attribute INIT_03 of inst : label is "556D7556BAAB7BAEF572CCBEB2D1C12D360037F4774AA01283DD2CEF6D12DD9F";
    attribute INIT_04 of inst : label is "9D3963451F7D948960016A9A84891C3A467C544500294B0A47A42CFAA64E4E5D";
    attribute INIT_05 of inst : label is "A86CAF17E3CB76DB6E3525D097247CE2C83CB7126F6A8BF29E6534DA693F95A6";
    attribute INIT_06 of inst : label is "92D209842B0517F44C91C3B9A81BAEBA29FEB534BA88D79773BE965788B2C922";
    attribute INIT_07 of inst : label is "9DDCF9E7F99C05E66D7594D6D4D67B536B1942DC90A01501A36448958FCD378D";
    attribute INIT_08 of inst : label is "804E4ED63127D995A0F76B3336C6E5A26FDC162DE2DE1631F7EC7DDC08E280B3";
    attribute INIT_09 of inst : label is "1BE4415CCB0364B113F55822224916F912602DF1C3431F20A6602DB258892D09";
    attribute INIT_0A of inst : label is "662DD5B25B2549A1C3BEA6AAB79E3C8F200825A0B5259BB3D3587F93B57C2860";
    attribute INIT_0B of inst : label is "CAD89FE7EA4F84EA0332E3BB28CF1118BB20AF6976952CF319A3F007D301C962";
    attribute INIT_0C of inst : label is "2606D6033B3333512E54976952E540134101A869B1A4836D2B5263023B1B5318";
    attribute INIT_0D of inst : label is "E0319733B137632FF960C130ADDBB02020211A82A01AD35AD1218D000BB3BB70";
    attribute INIT_0E of inst : label is "2035B7C0B26924CF678DF3004B6A1FF887B802B0C184A1229BE334D694B2B68A";
    attribute INIT_0F of inst : label is "1530AA67762E6B92EEBBECE4B143BDE991E446B98E11DEF6FB5B129A32F20809";
    attribute INIT_10 of inst : label is "64A73ACCE37127253519CAE24599C91292CCCE44A6ED99D91292CCCE44A6E666";
    attribute INIT_11 of inst : label is "6B1CF2ABA4B68197FDCA5B6F7206013C3A9ACC5048D96B0329242D06E7749862";
    attribute INIT_12 of inst : label is "DE703A0266FC5B0B4FFC96DBEA117BEF28957957EBA9A80BB6DE006F0641AA31";
    attribute INIT_13 of inst : label is "8136440E9287C6FB6FE07F1EB64441C2A9E1BCF9F3B0DFF5BB6DF5541007FFFC";
    attribute INIT_14 of inst : label is "C3E1FCF7E618BC01CB68FA8C723CA02BEB7FF0058804AB15145A0401DB64D3FC";
    attribute INIT_15 of inst : label is "64A910E1803FF6FEFBD9728D362AC8088A47303BBAC1BF8649380573A9027B97";
    attribute INIT_16 of inst : label is "FE88F9CD053A91E092422770E262DEC60395037B2E51940C54B5C0C0000DB6ED";
    attribute INIT_17 of inst : label is "D1750B68AB4F83EAD6430F4C849F3535D52C47504FB004FF47FDEEFFDA6CED96";
    attribute INIT_18 of inst : label is "A0CFF395F8DE5F2900136BD39C4FA2E0408C0B183A303B756063A1CA3941CE16";
    attribute INIT_19 of inst : label is "548050138E6BAA3BFBC7CE6829CA9B00138888897EF7FFB9FC4F78F7EBEB7DBF";
    attribute INIT_1A of inst : label is "D03FFAAA36901A9E7E0400670DE2CFF71F9268228A26E9FEF35137151CCCD444";
    attribute INIT_1B of inst : label is "C97232749AA883ABEC0CCB6925E18E0128073A9C1DB00E790200100A7F0BA046";
    attribute INIT_1C of inst : label is "4729F67BDDF080190498A4D5401AF26B3EB291049600099306490EF01BDACE34";
    attribute INIT_1D of inst : label is "E9234133801C03000599B588EEB3B3810454B1041094B67C92D2CC03319B7329";
    attribute INIT_1E of inst : label is "0EB63EDC4681D689E5B82B33F4B0C0D924F689B79300321072F24593B9D927BE";
    attribute INIT_1F of inst : label is "958392DA408040000586608000043FD88198C0601A00EABF12483800B03880E1";
    attribute INIT_20 of inst : label is "60602820004810200000200000006078783020105E689684EC64233F28D16A23";
    attribute INIT_21 of inst : label is "FFFFFFF951515151515151504151515151515151515150606060102008606010";
    attribute INIT_22 of inst : label is "0000000000000000000006606020001F01F080261305750301B4000404000007";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "6DB6DB6D6C89A9C766603F9FFFDF963C7F70210EE571EB06259C9FEF2BDD8DE0";
    attribute INIT_25 of inst : label is "04B5A0425ABC002BC3F9FC7C0B40B49C16EECA90599CA91FCFE5B2F98B05B6DB";
    attribute INIT_26 of inst : label is "427A9BFBCA1691688F1FCFE7F23E05A04B520521D7E78CA168F1FCFE7F23E052";
    attribute INIT_27 of inst : label is "6921AFB16265DBB936CB1FB82A2DC0A43653337831117F785152424A3C1D7F0F";
    attribute INIT_28 of inst : label is "BDD7FFFF5FC93AFFC7FFFFFFFDF3FFDEFFC05DD6E05DD6E0F0E69734FF8E7FE7";
    attribute INIT_29 of inst : label is "4810C0814308A38184410441044110002FF0FA82F8CD87F0F7F0FF83FCFE347D";
    attribute INIT_2A of inst : label is "BD60A343040A200088A428AAA230633332188C606264C088C649555555514444";
    attribute INIT_2B of inst : label is "A18E180CCC82306302360400C94BD303F4C0FC652F194BC652F1E0D7570C6EEB";
    attribute INIT_2C of inst : label is "000000000000000000EC262A16F1B77638D6C7D0F853EE5147027200000061B9";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "6E4A52A50FFEA6ECEE8FFE3DFE00EF7275770770757EF936761231272F4D85D4";
    attribute INIT_31 of inst : label is "6551503F0ECEE3F3CEE0EAE4C0DC0888990DDC13CEEEAEE0FEEE8FFFF0EEAEE1";
    attribute INIT_32 of inst : label is "F02DE60B1FCFFFEF1E2CEE2CE6ACEEEE0066600011660AAAAA4EEAEC3DFEE2F4";
    attribute INIT_33 of inst : label is "D2A79CA50A6CEEEEE8EE2AA2A2A9ABE7E0EEECEE6E88AA2E4466577737671990";
    attribute INIT_34 of inst : label is "000000002FFEE6ECEECFFF7FFF39EF7375775770FFFEF9BFFFDFFDFFFFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "087099CCD95EE30950E007001C0430100100100100104401C3C1593693113000";
    attribute INIT_39 of inst : label is "7837C17CBF33C4BE7E666C978565DBE7913102004126CF024D9A01E00700C593";
    attribute INIT_3A of inst : label is "18020000C0189111ABEF94905933E7B3ADD9F92ECFE4000DE001ACB2F0017216";
    attribute INIT_3B of inst : label is "FF812250205305313A2C0263B924B95BF2504A0201A8792B00C1AC3C94BE0522";
    attribute INIT_3C of inst : label is "192F4C93A65876192F0C978649C324E192F0C97A64804100BFFFFF024504804B";
    attribute INIT_3D of inst : label is "023804C03C01FF80010C80406DD41880618649C324E192F0CBC325F8649C324E";
    attribute INIT_3E of inst : label is "000000000000000000000000000000000000000000000000000049B36DED0189";
    attribute INIT_3F of inst : label is "1200000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "76D86BEB05E860CE1F522A83070E24550A04301982AAD4006E00000000000420";
    attribute INIT_01 of inst : label is "81FF0397E676DA5152377FF70FE5C8E168373923EC70859AC6D93FC2E37D9F5B";
    attribute INIT_02 of inst : label is "491B4A366A93350E6EC22AA5365F6B2FB426997FAEDDCA9AEDC37E2946824D1F";
    attribute INIT_03 of inst : label is "CA0A022F755F555112C087279CBD4DB99D28E87EDA7B484AA003FDB44D909DDA";
    attribute INIT_04 of inst : label is "910FE2034E7C8C1796C7BEEDA6E8148B444428280508428AAD21005046464671";
    attribute INIT_05 of inst : label is "B9DC1F23F0026DB6D475205953022530071C0D986F5C800213042E085B1FA945";
    attribute INIT_06 of inst : label is "2E2B085928DD2F5400086403E15A32020980FB9CC5FE1D188BB1FB54ECFF6D33";
    attribute INIT_07 of inst : label is "354550260005922B091F3984798478E63F12D48C0384B450852A408BDC3D2C59";
    attribute INIT_08 of inst : label is "22040221A401B00AA830358126728C7A28987478E78E3A2054C21545811A805E";
    attribute INIT_09 of inst : label is "7B57366F7DE7FFD9B5E67FBBBB583C50B61478A1659DCA9B37BCF7FFECDA4B1D";
    attribute INIT_0A of inst : label is "7F7677FFEDB604A0440B9D959070FC3F103DA9282B03385959D46000800D6034";
    attribute INIT_0B of inst : label is "571E76FDBFA1069BEDA092DA4A49B9D9BFF56C7E5BE5B7ADACB9A11002092833";
    attribute INIT_0C of inst : label is "DFBBE134C81BB9792B6EE7FE7F10A86DCB4B72BB5829155779BAD75715CEF401";
    attribute INIT_0D of inst : label is "F13EAA522912139FB15C9558D1A23001381D1C8B200740E82EEEC3CC689B3179";
    attribute INIT_0E of inst : label is "050031D402B800525527AD884DAAD7E90FEC31AAA128397F6ED22BF7BDB6B2CA";
    attribute INIT_0F of inst : label is "C9964A4554368CAB6ACA021C0042DE4A80C220B0EC916F32A10904B540375B5B";
    attribute INIT_10 of inst : label is "4AE43EE83A2AB05729106C55604242A0842152A820884252A0842152A8209772";
    attribute INIT_11 of inst : label is "B8FC7149740AA152D5C55601750495112B5CB61C440A5502055603D445DC95B0";
    attribute INIT_12 of inst : label is "BE5C337EA155C5E1925D1410F31DBAFEAD1F61E6292815BBFB6F6C346301701A";
    attribute INIT_13 of inst : label is "3F001C4A850554D250408B97B50001C21172808102B91925BFB6E9A7D01544F4";
    attribute INIT_14 of inst : label is "AFD7F421615AA3C16DAC7AC755C7ED83E987A6C1DC46D7AA5D78B2417E3E0680";
    attribute INIT_15 of inst : label is "5FEDCEBF88A528C84830438E043F6C448A8538272A5D12A54102512150055237";
    attribute INIT_16 of inst : label is "960468E94B0B9D38A17ADE4833BC736F7C46A3B60871F96A7EDD628A408B7FB6";
    attribute INIT_17 of inst : label is "D1FFFA68FDBDC2AA16D5A7C1E5F9DEFDF7EC48504D2204A5840E634C824F89A2";
    attribute INIT_18 of inst : label is "3E8C00AD7ABA334795FD0880CE9557F0478CC86910D2FA220073E1FA3F59FFF4";
    attribute INIT_19 of inst : label is "642ADC3CEBFBEF5203A3474A584B1E21031D0D12C0425285F4E614A14EF84620";
    attribute INIT_1A of inst : label is "D21B680A1D0EC284428D4A6361C28C065971E71E785C4180DDDDDDD997677766";
    attribute INIT_1B of inst : label is "F9217058CCF0892B5C87B1BE374384443AC755ED4DB2ADA11712B61311E0A413";
    attribute INIT_1C of inst : label is "67E9141F9BF4EDD2B6D5285D68106351143480011988C914246A2A191E186F90";
    attribute INIT_1D of inst : label is "8809D016A455224BE000244020242219000448AFECD902951B50B90229580B2D";
    attribute INIT_1E of inst : label is "08B39458ACDC8002CF900B59F689A2FFCE800FF939885A38A0342000D0FF5A9F";
    attribute INIT_1F of inst : label is "AABFB4D830800000070879010002503E81E0858269006077E484150040010001";
    attribute INIT_20 of inst : label is "1010181078304010303050303030107878781058178CF33D762C0DA266066F19";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000101010401038101040";
    attribute INIT_22 of inst : label is "000000000000000000000878402000AAAAAA02000305751303B4040000000800";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "1208208241492B554A6BCD274E9D25695541940B494B5A4203E94A5A4969487E";
    attribute INIT_25 of inst : label is "18A2033120C93642A2A5509065225012648A9108921D10152A8104D52A020104";
    attribute INIT_26 of inst : label is "99D2955692CA024852550A9543C812018A213286955A492CA52552A854BC9129";
    attribute INIT_27 of inst : label is "FA01691912445092269255240A0D26522092A2D21114AAD128404049696954B4";
    attribute INIT_28 of inst : label is "42085540095990C82509011005092AA72AA309054348014338482A2555571553";
    attribute INIT_29 of inst : label is "004440ABAD8880C010541054105418010FFC8215550890500250014040A02052";
    attribute INIT_2A of inst : label is "42C5543E245577FFDD6B77FFF76140010000020C401C600020B0AAAAAAB06000";
    attribute INIT_2B of inst : label is "9D7DD620154C4C84CC4C151982A5ECF92B3E4A8A97A2A5E8A97A438A8AF85045";
    attribute INIT_2C of inst : label is "00000000000000000016F1B77238D6C3D0F852EE5147FBBBFC0944BBBBBBC60A";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "D423F3EE09989198BB8BBA3DFE11899880880FF0B026603EEECEECEF2F4D85D4";
    attribute INIT_31 of inst : label is "D40D74550B9981910770BBA1B2B82EEAFF0BBA13033330101010000000450DC1";
    attribute INIT_32 of inst : label is "DE6F6C50130111091A39AB1DF7BCFFFF11EE7BF2FBEF1776775763743DDCC0D4";
    attribute INIT_33 of inst : label is "F206B07C0A311111107F6737F7ADEFE7E0777477321DD80D5DFEDCCC8CCD5DD0";
    attribute INIT_34 of inst : label is "000000002FFEF7FDFFCFFF7FFF39EFFBB9BB1FF0BEEEF9BFFFDFFDFFFFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "5211C088004FF0125AA01501128E1A38830830830A38401453C0F2DB6C881FF2";
    attribute INIT_39 of inst : label is "FC085BB49E000DDA3C062802DF790CEC8A70020D010A4F82149B03A915480D00";
    attribute INIT_3A of inst : label is "C958001348CA81311000000098536283C341F81A0FE0C9066C9067272648370C";
    attribute INIT_3B of inst : label is "AD280144C958158548C1586771B6FAD3F5615054AC0111C8561628C8E444190A";
    attribute INIT_3C of inst : label is "925E492B2492449256492B2497924BC925E492F249FFBEDBEAD55A5003DFFFB6";
    attribute INIT_3D of inst : label is "820B25605520407FC1EA846D099C1280412415924AC9256492920AD2497924BC";
    attribute INIT_3E of inst : label is "000000000000000000000000000000000000000000000000000042934A8A42A9";
    attribute INIT_3F of inst : label is "7C00000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "56CA20F345AD56760F0ABAD96B0E1574B4CD90010A6992003500000000000044";
    attribute INIT_01 of inst : label is "8150439784E8F0AFAA6D77A146C1C8F478989FFD1D109D9B4B6BA4CBC7A4D951";
    attribute INIT_02 of inst : label is "025F587DD1DEE8A726A82AAF9ED5256A926AC8699659DAB2C969682242C34A2C";
    attribute INIT_03 of inst : label is "4AC3EAC8656695D56280ED073438F594950A81C139174A0261AE4272A3C70313";
    attribute INIT_04 of inst : label is "C437A37CC2ACF0C49255AC2D0653C5B1C38ABEEF050D088E48061167C1F351C5";
    attribute INIT_05 of inst : label is "150681B5B0827FFFFC452489F10210D419588910187E8402918D23585953D09E";
    attribute INIT_06 of inst : label is "BA7A20F1E9713A1404084283C04C90820D34CC8DE665CB1AB2E6495155492599";
    attribute INIT_07 of inst : label is "A3BB8034D0849E1EE11FBFC47F8E53FE3D1B98C40320110621840E1F59DCA1F5";
    attribute INIT_08 of inst : label is "C2060237D901F83F921E3D86598E0FFC5188C378D7C23E341A8B05AD8409C1E8";
    attribute INIT_09 of inst : label is "4C7B122AA4F49248F4FAE799997FBE402FC57C805ADA8389155E924924794706";
    attribute INIT_0A of inst : label is "555ABA4924920448570BB3BBA39630AC237F9C102B045F5838E14D008106425D";
    attribute INIT_0B of inst : label is "8ABCF23C8EDE55B6FE2DB8D51F288CCBFFDF663A2FA2F3858E3A35581BA48191";
    attribute INIT_0C of inst : label is "DB7D764FF3135B98A7B5A2FA2FC11824CB6B12B9DB449677198A7A51BDCE3334";
    attribute INIT_0D of inst : label is "75503FC57E39F99D71E2E2704817681059231589CAA69CD336972DDBF3935B9F";
    attribute INIT_0E of inst : label is "757D26D5BBF16951F2C305A8C2445AE1C8460B9250C0B8790E63FEF73D8E7BAB";
    attribute INIT_0F of inst : label is "CD96ECAEBF66FEB66FEBC268A0CBBE53DF8AF4EA597DDF3CFB7E149E74B45B5A";
    attribute INIT_10 of inst : label is "265174A55A399132870AA063204840911424522445C04840911424522445DEF2";
    attribute INIT_11 of inst : label is "E4B8A37520DCE2CC9C8D6C60BB8B1D1E099456C3158D1A89043344E0600A4A37";
    attribute INIT_12 of inst : label is "C272016001114711B0E6C1C7BA0041873970FB0EAD6114947FF127351362A39D";
    attribute INIT_13 of inst : label is "442BBE9E1329A9C83030EE3C13AFFE6038E0AAB52A30409B47FF018E23326909";
    attribute INIT_14 of inst : label is "DF6FA894C5700C104240F909760B64D9049812547852FDAAD9689CC6DF6E44D6";
    attribute INIT_15 of inst : label is "12F7E5342AD60C6C75A6FF0747F32D51642334158842684D4E3806C485838DB2";
    attribute INIT_16 of inst : label is "62BBB170830D699C316C4C5811157B695702E0B4DFE0FBCFE6C86BDE45864BDE";
    attribute INIT_17 of inst : label is "EF9AB0F7CDB0E1621C61613DE1E017BEEBC46887669AB4722DAB3DCA4A09413B";
    attribute INIT_18 of inst : label is "3F69A08E2C2C47FF857B51109DFEE8182F4FB1F7B3EFD2627051E8ED1CA0ED61";
    attribute INIT_19 of inst : label is "21C8DCBC897DD798D21D8B841879B4A8510A5E2F984A52CC831CC520407F0A8D";
    attribute INIT_1A of inst : label is "EAE80A8529D4C3667285025522F069A589AA8AA8A3778D348C8CC8C8A2322232";
    attribute INIT_1B of inst : label is "F92FFF9E6C312D374D8A92F25E6B60243403112889184622CA091D13071855F0";
    attribute INIT_1C of inst : label is "74CBAA65B940E4B7D67E16DC6A90F3F559DF15842E0A28120111A35B178E6F9F";
    attribute INIT_1D of inst : label is "91B81014A444058F5C1C38E8E424AB515418CD4F6A5D6B02CBA3F9537C4788AC";
    attribute INIT_1E of inst : label is "854C75407A829012AF08C6A7B0F0EEFEAF20076DAAAAEC12A09485049CEDFD75";
    attribute INIT_1F of inst : label is "C0E380688887F800050000000003900A19FD821A04004033001016FC40165441";
    attribute INIT_20 of inst : label is "CCCCC0CDA2A0EFCFEFE8CFEBEDE8CD828580CA8287F29220400805EA2A00324D";
    attribute INIT_21 of inst : label is "00A2000000000000000000000000000000000000000000C8C8C8ECCDE0C8C8E8";
    attribute INIT_22 of inst : label is "000000000000000000000F8321800071C71C0400032577032598000000000002";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "A4D34D3448490C62363181D16045D32E6EFADDBD34B8178003BEA423A4ACD460";
    attribute INIT_25 of inst : label is "285BB7B24C867BE3A379BE3EB64F66FCA76E6D939D9AD9BBCDF0A0BFC584DA69";
    attribute INIT_26 of inst : label is "6D5C1FBBC36CD84E819BEDE6F89F7B3285BA7B3266EF8836C839BCDF6F09E7B2";
    attribute INIT_27 of inst : label is "B76129557AD5FB0DA46D9BF8090BCF74A4175F5CD5D9FD7FB333733A262E6F1F";
    attribute INIT_28 of inst : label is "5E6C7FC24B7038ADE3F6034F05E53FE53FF55D54F51D54F528E287A57FD55FFB";
    attribute INIT_29 of inst : label is "145100C10408800540554055405540250EA279481CECC7DAF2DAE3EBBEFF347A";
    attribute INIT_2A of inst : label is "0002002802080888008020888003400455C00106400048001000000000010000";
    attribute INIT_2B of inst : label is "8828811555550150150055400004155405550000100004000100060888A09440";
    attribute INIT_2C of inst : label is "0000000000000000007238D6C7D0F857EE5147FBBBFC1510540011000000028A";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "386846A1077EF770774664044411EE2471FF0FF0B895F818991111190D4F86E4";
    attribute INIT_31 of inst : label is "12E53A38071767F78FF0F761F6FD3333330FFE118FFF3CF2F6F7B7D7F3FF2FE3";
    attribute INIT_32 of inst : label is "B06D2EF50E0FEE6F1E7DCD1BB330BFDD11CC59D0C8CD1776775763743FFCE2F4";
    attribute INIT_33 of inst : label is "114701950E79EE6EE87F6EAEF7AD666760DDDCFF3E5DD80D5576667717667FF0";
    attribute INIT_34 of inst : label is "00000000277EF775774FFF777731EEEEFDFF1FF0BABFF99DDD9999999DCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "1A11C0B4C04DF4007A2911003824A29A09229A29A29AAC144181FFEDBE88150E";
    attribute INIT_39 of inst : label is "EE478B889F13E5C43E24148E584ABADEB16803650060C9D0C193822911003A90";
    attribute INIT_3A of inst : label is "59030050281A1111E8000002091924F16278D9138406881D68130966B409B311";
    attribute INIT_3B of inst : label is "086002A0450350243945033B34925192F3150A52818295094088390AA4A50128";
    attribute INIT_3C of inst : label is "2BF79DFACA6CAB39F594FBCE7DE53EF39F794FBCE7FFFFFF55B810D206DFFFFC";
    attribute INIT_3D of inst : label is "D06A25F064004000192AB40C0BCC2A8062CEFF677EB2BF79DDE57EECAFDE77EB";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000000000000000000000009832FF5598A9";
    attribute INIT_3F of inst : label is "B200000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "564A61C340A47446C05890095360B1201050120204D22410F1020000000000CC";
    attribute INIT_01 of inst : label is "125A4421757C589A2BB721274DC1CA64397CFDB30C3891CAD6596D892EADDB50";
    attribute INIT_02 of inst : label is "681882B5435BA1AA6CE02AA987740EBA06D2DC79A6DDC894D59B682948594832";
    attribute INIT_03 of inst : label is "86414640A3200CA32AE2D463D1984C9CFC088B405C031029233A00B881C28281";
    attribute INIT_04 of inst : label is "003A06286A2CA08DB6C58F8E26C14191D0982241552C09AA45050B230545E751";
    attribute INIT_05 of inst : label is "3148C81AA24976DB6E944661172640E24C2CB5209031069E8895172A35506945";
    attribute INIT_06 of inst : label is "A0A0C1432A43A350DC994AF4054A02126D129998ECCC1D119A22DB56EEDB6D33";
    attribute INIT_07 of inst : label is "345554D4499668E10D69A0CEA0864183503B46DC9486844283A40C1C68E870C3";
    attribute INIT_08 of inst : label is "2CCA4A828525D898A810DA130F4A0C4841C147C81CC06067549FD5100EE15132";
    attribute INIT_09 of inst : label is "4526B6F67F8DB6DDF806B7BBBBC0E6023807CC05B9D9895B7BB1FEDB6EF00024";
    attribute INIT_0A of inst : label is "BBB766DB6DB6CEC0851419110353D1D467112B28A7255A2D1D45449285D9833C";
    attribute INIT_0B of inst : label is "1D39CA328E4D589C644C98C87C23B9AFE89AD7B09B8DBE1FB03411100002E177";
    attribute INIT_0C of inst : label is "7B4D644AA3F7DD98A12009B8DB50996D95947D3D180C6A4771BF4DA7318EFA80";
    attribute INIT_0D of inst : label is "311FC2499431210985481062532233121219148B289AD75AC39309936377DD9E";
    attribute INIT_0E of inst : label is "1A04A3281D410484412E1F8925A30A009E2425B2E42A4313C6432B435DC6075C";
    attribute INIT_0F of inst : label is "29594A45015E569DE7694660A0C26BE122444292445935E8508411D30058ACAC";
    attribute INIT_10 of inst : label is "2D145CA9923B4968A913287691DB6BB6BCEDB2ED8CB9DB7BB6B8EDA2ED8CAEEB";
    attribute INIT_11 of inst : label is "0768A284E0A8655A888A14F7B694B91821149C8B5D89540A30684B64644850E4";
    attribute INIT_12 of inst : label is "C364903FAE01F84F12C11410B444B90100D27537C0A1D5B65B616F63962507B3";
    attribute INIT_13 of inst : label is "32631E0836A0E5DD60659A059600000B7504A081422240CA65B61DFE9ABB320F";
    attribute INIT_14 of inst : label is "B25934A94478068524818718234FCDC305CC16D3BF66D52A596895CB7CBE944F";
    attribute INIT_15 of inst : label is "46CDBC7408E7878C62464E1644E3B458AA84792E090822A6482E4080502C7310";
    attribute INIT_16 of inst : label is "823401894D29F1003A28DC48F330716E55446738C9C2D209C76CE27E4B9D1B37";
    attribute INIT_17 of inst : label is "F7188CFB8E6DE68E501235100F4C8ED065A35014E8248CA42C92214C186E8D83";
    attribute INIT_18 of inst : label is "B22892B56A80731271A001328E154899688E018C1719322ED0D2894328614119";
    attribute INIT_19 of inst : label is "60AAA18A49A0CB684BA00C4A69513440C328284909C631D8075EDE6D38181A84";
    attribute INIT_1A of inst : label is "424348D824587A367B02024CBCA4209645C71C71C64F1D129D9DD999A7766766";
    attribute INIT_1B of inst : label is "76C4C41CE47408E73F9AC5B8B6234506820422945068214805102AA5E5AD849B";
    attribute INIT_1C of inst : label is "6AE176E2AD30ED823245AC58703963124894108D59504C12810140272E2E439D";
    attribute INIT_1D of inst : label is "814D032A8894404A61CF31904DB223E108B0E809B0DD24D19B023206090A382C";
    attribute INIT_1E of inst : label is "287A5544618860802672C5958080D644A7709EDED98FD85892800092CA26CAD9";
    attribute INIT_1F of inst : label is "2F100602277800000287FB83806420503DFD4449138088C4E6CF000015000014";
    attribute INIT_20 of inst : label is "A3A3A7A4A1A780A0A0A7A0A0A4A7A3818487A6A1A7F265888641A05100C1005A";
    attribute INIT_21 of inst : label is "288A8AA820088028880088000008A0A008A0A8A0000887A7A7A783A4A7A7A787";
    attribute INIT_22 of inst : label is "000000000000000000000FF8000000FFFFFF403FC74575030200404040404040";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "5B2CB2CB6DCE46514E29243408953401510026000D6026466789884A65290CF4";
    attribute INIT_25 of inst : label is "0034424D32A9201A4685404009A0984204C01A680311A20522843691242B2596";
    attribute INIT_26 of inst : label is "C21213401A130B694A540A1501200440034D24C295084DA114A542A05092104D";
    attribute INIT_27 of inst : label is "920DA5512B849103349854042929249A36DEEC021994620049AC2C6501295090";
    attribute INIT_28 of inst : label is "E4D7D55F38C806B6550D04FF5502EAB9EAA261B22261B222CB0D9135D5597558";
    attribute INIT_29 of inst : label is "E0A2000104063E0ABFAABFAABFAA800460808305510BC8390E3914A440802E4F";
    attribute INIT_2A of inst : label is "820444382022AAAAAA2A8A222A8140020740820C42086008208199B9B98306EE";
    attribute INIT_2B of inst : label is "88288008000800800800AA8005D08020200809574255D0957425068A8AA0D4C0";
    attribute INIT_2C of inst : label is "000000000000000000C7D0F853EE5147FBBBFD15105440545404444444440282";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "902FEC4488088198BB0BB9BBBA11EF3CD9FF0FF4FEB5F838AA2EE66E2E4707F4";
    attribute INIT_31 of inst : label is "BC516ED58E8080808880C4C0C4CCEEE2EECEEE028CCC0CF0D4C484C4C0880983";
    attribute INIT_32 of inst : label is "143F94410F1101191C5DEE0EC9D49DCE22CC7BF242631BBAB39BAAA82AB02230";
    attribute INIT_33 of inst : label is "B902EF040C510111101919988088088888ABB8BB3E3BB80BBBFF7EFF9FFE6FF0";
    attribute INIT_34 of inst : label is "00000000AA2ABBB9FF4FFFFFFFB1FFFCDDFF1FF4FEBFF9BFFFBFFFFFBFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "CA510960C95CE00974A225107D30E4C34C34C36CB6CBB554804189A6D31925A5";
    attribute INIT_39 of inst : label is "447FA18C0133D0C602622093A407A95F3D0983B481EBED83D7DB04A225103413";
    attribute INIT_3A of inst : label is "32060048923A117BA8000000413806F36571812B8C050A14B03300AA6818AB05";
    attribute INIT_3B of inst : label is "054D031C0A07206022260704C124A1500242061303A0712981D1007894880530";
    attribute INIT_3C of inst : label is "936649B720C204836E49B724DB106D8836E49B724D34D34D20540A9A0749A69A";
    attribute INIT_3D of inst : label is "82CC04E0B4437FFFFC402919C9EE14080120DB906CC9366498906CC20D9106CC";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000000000000000000000007AFB48887ADD";
    attribute INIT_3F of inst : label is "B400000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "A490429A49A5A2DE4869080B3F20D2101EC5BA0B5E9E7402740200000000048C";
    attribute INIT_01 of inst : label is "5BE909582562010C2BAD200209557F406225A49009268D3C9413297BC72900A6";
    attribute INIT_02 of inst : label is "446492B4591A2CDF6FC9D7E1855545AAA23BD54DF69DC084C3793864AA794B60";
    attribute INIT_03 of inst : label is "E6592ED2B3211DA3278AD55A55567DBFFC9B080990125884086053209176A8AB";
    attribute INIT_04 of inst : label is "56A840C45EFC91ADB6CCAC2D926B5DB766C8C8AD9BAC6DAAE76D9B66155555D3";
    attribute INIT_05 of inst : label is "2669A8D85A5940000BD40D421376D5A7587EAAB7B02332634846908D35D47B6D";
    attribute INIT_06 of inst : label is "50D081A4BBA4C7F2DEBB4A8E80FA42DF6E92D553AAA911519DF2926088924966";
    attribute INIT_07 of inst : label is "7CCCF27E4BD400672D70C061806B6300C20506CEDF8075D8B68F6AD4A48685A4";
    attribute INIT_08 of inst : label is "35EF5A6AC7AD06B0AD3261577E0A1C86D97017031064049CA28B290EED050212";
    attribute INIT_09 of inst : label is "842424554909249500255F6EAAC1838040490701C53F21122AA124924A8B6C46";
    attribute INIT_0A of inst : label is "AAA5449249246D85D938515556121084264925AEA76F793B1B43E4D6972C0620";
    attribute INIT_0B of inst : label is "DE19C22088D44592DD2596CC7961112BA800F7BACA28342938A11727D5010B22";
    attribute INIT_0C of inst : label is "722E4D20895557138258AC328356824954152521536DEAD425145EA2752842B5";
    attribute INIT_0D of inst : label is "26FE92C60B6A1FEB03259DBB7B768520BB344E2FACC895125B8B9949F9555715";
    attribute INIT_0E of inst : label is "6A2CB2E9BC0B65DC1734A9307818490093ACA657E9399583265AE04217CF0E3C";
    attribute INIT_0F of inst : label is "29414B98CD0EC2B0EC2B4EC59256395B4402A28200531CA2D4A5371776E2A0A1";
    attribute INIT_10 of inst : label is "A2832D6498B0A5141189256140C949921064C26487A8C959921064C26487B768";
    attribute INIT_11 of inst : label is "8D14F29CED9008954E4A0869312204DA9FAE60600CE92029AA14241373584C02";
    attribute INIT_12 of inst : label is "C5E117826A0E2B293D80B514E74F03A18E10E50E40EB292AE921DB0010C8C280";
    attribute INIT_13 of inst : label is "4426261811B4C34810232934B1401F4764B563C78F1AE08EAE920BAF1230200B";
    attribute INIT_14 of inst : label is "C2E162C215DB6E4CF818C18D33ADA908050816C40D96FCDFDB61E61258AC484C";
    attribute INIT_15 of inst : label is "82A549AC3904A65DE1B0CA252CA249A64BB6BA377C656BB05B7ADDD6774A7351";
    attribute INIT_16 of inst : label is "5AD48B4D676B8B5A727896C1AAA55270B95A08361944809944974448D0A40394";
    attribute INIT_17 of inst : label is "451024A2892B4BFED119AF0E55084C10416CD8C41EB601F6BC9A657A19684D0B";
    attribute INIT_18 of inst : label is "EB3C969FFB42C32158909B16AE4516B291AC7B18523022A6653A894128294049";
    attribute INIT_19 of inst : label is "5D994AC02820827E4EA45A6B3B5FAD6128AAAAA08CE77985821C4C2E38994AE4";
    attribute INIT_1A of inst : label is "C0217BB8C2A9420F47B30D51604934946D000000018C4F92DDDD955557755775";
    attribute INIT_1B of inst : label is "524C4CD6A1AE30E338A0D432942714D5837000800030010001C002B9092B8056";
    attribute INIT_1C of inst : label is "57EB20E6A9222956B489ED5358054A2759B2B336C2980C57D01B64384BAFC2FB";
    attribute INIT_1D of inst : label is "EB2B0FBE81D40872A5DCA14ACCB96A350515844490976ED59216430091291AA9";
    attribute INIT_1E of inst : label is "4DF05DC6D26472DBF51A5D05C19F9E403502CA90513210B31676CDD2CBFF121B";
    attribute INIT_1F of inst : label is "000600000FFFF80000000080806200003C004000000000000000801154801154";
    attribute INIT_20 of inst : label is "202020242720202020202020242027070300210000048000030180600400000C";
    attribute INIT_21 of inst : label is "DF5D5FF82028A880080880000008A8A0A8888080880080202020202420202020";
    attribute INIT_22 of inst : label is "000000000000000000000007FFFFFFFFFFFF1000230775230000404040404047";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "4B6D92D9B6EECED88DEE4D370E1834E9D5CE4CDA0D666277F7C9C3526D692EF2";
    attribute INIT_25 of inst : label is "A2B98C9092E1C98A22A351D1921D31918CD91CC73355CC551A8B5AC2384925B2";
    attribute INIT_26 of inst : label is "64D3D356AB2475AC3A751A9D4F69E99A2B99C90C9D5236B263A751A8D4768E98";
    attribute INIT_27 of inst : label is "F662B5156255B393559A7526A8AB39235B5888D355566AD68E119891E1C9D464";
    attribute INIT_28 of inst : label is "433055609CDCC2C83D1BF890FB192AA32AAE869B2E869B2E1C34D956D56BB557";
    attribute INIT_29 of inst : label is "40F300D6581EEE0FFFFFFFFFFFFFC016E9958AAFFBA9813027303C40C5A2A54A";
    attribute INIT_2A of inst : label is "D706EE90201101111100544444023757529DD75B375D3DDD75C199B9B9830444";
    attribute INIT_2B of inst : label is "2382281DDD5D55D55D50FFC00080802020080802020080802020042020008195";
    attribute INIT_2C of inst : label is "00000000000000000053EE5147FBBBFC15105540545411150100000000000131";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "AA8000008F7FE6E8EE0DD9FBFE11CF3CFBFF0FF4FEB5F83DFC1DD55D180B8194";
    attribute INIT_31 of inst : label is "AAAA80008F97E7F78FF2F383F4FDDDC1FFCDDD17177738B0B3B3B383B3777743";
    attribute INIT_32 of inst : label is "AA8000000F1FEFFF3813771FCBF4338B33883BBB8BFB1DDCD5DDC9DD58D5FFF0";
    attribute INIT_33 of inst : label is "AAA800000EFBEFEEE0FF7FFFF7AF7FFFD9CCCC444C22200999DD189B999B2AB0";
    attribute INIT_34 of inst : label is "00000000FF7FFFF9FF4FFFFFFFB1DFFCFFFF1FF4FEBFF9BFFFBFFFFFBFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "6F512DF2ED4DD6ED66A075026D30E4C34C34C34C34C3E66ECAED8DB4D25DBE95";
    attribute INIT_39 of inst : label is "54F7DE8B81A7EF47034832D2F486897E6BCD072F8B369B066D320FA07502265B";
    attribute INIT_3A of inst : label is "1F03800018159B5DA80000005D335538629C2514E1158064B80610AA6C02AB41";
    attribute INIT_3B of inst : label is "FFE08A000302B03B2027038001B6E9D5034B03B381405529C0A0002A94952538";
    attribute INIT_3C of inst : label is "D16668B730434CC16C60B6305B1A2DCD16E68B7345A4DA4DBFFFFFC1164D26D3";
    attribute INIT_3D of inst : label is "07D80E41D40F7FFFFD000C0F2B8CDE1315305B982C8C16660A1A2C934599A2CC";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000000000000000000000004DA64A984D83";
    attribute INIT_3F of inst : label is "B800000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "76DB24C36CC94446994A3BD143429477A09D104D5A0C5000DE03000000000101";
    attribute INIT_01 of inst : label is "80FF79F18056795D6223BB7165C5C27628B5B24B0C98D18E4649AC89AD6D9B51";
    attribute INIT_02 of inst : label is "005659FC823E414C6D842AEDB4574A2BA4E3D97DA6DD9BB0CFCB78205682280D";
    attribute INIT_03 of inst : label is "0000089AD44D513452B047031C19C5B8150A85ECDBF36802A0ADD9B63980080A";
    attribute INIT_04 of inst : label is "310DC840CC5E806DB6C5AEEF06F0C401618694E3FF0140020D01105440C0C041";
    attribute INIT_05 of inst : label is "11929013708009249A640484E6000830030C1D12380F24808200040201144186";
    attribute INIT_06 of inst : label is "8808801478941D50040003860048981404A4088CAC44DC022994DB02665B6C11";
    attribute INIT_07 of inst : label is "044450129081922000061900990068644E00B4580B0020000122C18295141814";
    attribute INIT_08 of inst : label is "A2120081B500280749B084810E4204300010613513049C045051140444180058";
    attribute INIT_09 of inst : label is "514336332D8DB6D8A40379B333289884A217310834C68A9B1911B6DB6C500005";
    attribute INIT_0A of inst : label is "999622DB6DB684881583222220D4D515406D8048080238090901290005080214";
    attribute INIT_0B of inst : label is "05945AB6AFCF40B3CF04B0C310608898EDB9463E4BE4B6C58132A51C710E30B1";
    attribute INIT_0C of inst : label is "238466033211115C837FE4BE4B60486D824210B398000667108CED1139862780";
    attribute INIT_0D of inst : label is "35908A001802310B411FD730C1031F08701E2D175FCED1DA71010D8002111158";
    attribute INIT_0E of inst : label is "414505052990490631A645A8DA42D5097FAC3EB1FFA09F1C60223F7399C6061C";
    attribute INIT_0F of inst : label is "9C24E466678EA2A8EA2A601820433942BB2EE40CE2059CA48E76113B14841212";
    attribute INIT_10 of inst : label is "2E442C69303397722D9260672D121A24A2890A8928ED121A24A6891A8928F544";
    attribute INIT_11 of inst : label is "99F450E400082046C74306A123017098AF0CA28E114D4F0A0C7348C2755C5615";
    attribute INIT_12 of inst : label is "D47FD10203040EF982C874F37E1345A994546146041015BAE4916CB16BC07559";
    attribute INIT_13 of inst : label is "0D4A060E27A946D4705FED1EF70443BE1D60B8B16290009FAE490597EFF10908";
    attribute INIT_14 of inst : label is "8AC56814A01003DD5A414397559FCD91059416E05D02D48B1860FE415E2E8694";
    attribute INIT_15 of inst : label is "32E5843E0894CA2420E06286062B6D64C2003782081E06AB401806E181F95A11";
    attribute INIT_16 of inst : label is "26081060420591A67338DC5819BC7979FD8120BC0C50D8CC56D8620BC486CB96";
    attribute INIT_17 of inst : label is "515CEA28ACBD829A0010E6047C70C3DD75C42804090A00A0ED216089C0032063";
    attribute INIT_18 of inst : label is "46E520085A241B05D2DC40A00C2BF6B0920CC021144268288038FC7B8F7C79D4";
    attribute INIT_19 of inst : label is "2008CF8C61BAEB4890C08302103F6EA011080801C142529C864694C10A888189";
    attribute INIT_1A of inst : label is "C005C890892DC402C0A108C0604AE52340288288203994A44CCC8C8C93333333";
    attribute INIT_1B of inst : label is "724646186E342C1E0482B0BE1743707C80CFFEFFFFAFFDFFFD3FFBD717F90032";
    attribute INIT_1C of inst : label is "7761B6231884ED8356C52858684853149551070C4FE8E4108000A3410E0E0388";
    attribute INIT_1D of inst : label is "901910468064075BC00440C42110061101283B96CE5C48954B202D090C10842E";
    attribute INIT_1E of inst : label is "F87218C40A5EB090E29647114388B36DE380865948AE582AA0A0850456B72EDA";
    attribute INIT_1F of inst : label is "FFD9FFFFC0808007FFFFFF7F7F9DF87FC2027FEFFBFFFFFBFFFE014150001450";
    attribute INIT_20 of inst : label is "808087848787878787878787838780A0A0A780A0A0037FFFFAFE7E1FF3FFFFE3";
    attribute INIT_21 of inst : label is "0000000000088888808000000008A8A8A02020202828A8808087808480808780";
    attribute INIT_22 of inst : label is "000000000000000000000FFB61A1FFFFFFFF0100030D7DC7CFFB838383838380";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "8240209200096F576AE8B3A0E1C3A0152A6994ADE8409142413D1DEF439C085E";
    attribute INIT_25 of inst : label is "19A29321001536406150A8386402403A668CD1089A1510AAA5518029A1FA4804";
    attribute INIT_26 of inst : label is "992A10A9C0C84002454AA542A19C12819A28321152A7400C8454AA552A19C120";
    attribute INIT_27 of inst : label is "D348000140051A3A80D54AF40001A6528009992A111415392100080115152A8E";
    attribute INIT_28 of inst : label is "46182AC08840B04877890010518C1563157B00011B00011B180008802AC30AB2";
    attribute INIT_29 of inst : label is "40A200000001440AAAAAAAAAAAAA803C45DF426050088010021014C063702042";
    attribute INIT_2A of inst : label is "8204441020110111110054444400000202008208020820082081111111020444";
    attribute INIT_2B of inst : label is "00000008000800800800AA800AAAAAAAAAAAAAAAAAAAAAAAAAAA054545008080";
    attribute INIT_2C of inst : label is "00000000000000000047FBBBFC15105440545411150150511108888888880000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "000000000111011155066062662202202222022022313035743FE66E2E4B83B4";
    attribute INIT_31 of inst : label is "000000008D9181130550D1C1D4644440664666268EEE6CF0E4C404C4C0880A83";
    attribute INIT_32 of inst : label is "00000000091101111C59DD1DCBFCB7CD11883BB989DB3BB8B33322646220AAA0";
    attribute INIT_33 of inst : label is "000000000CD9898991555444440444CFD9EFFD7F7CBB7C4733753EDDDFDF3AB0";
    attribute INIT_34 of inst : label is "00000000555DDDD9FF4777777733D66477771BB02237313FFFBFFFFFBFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "4800C06C401B34000A201100010014004004004004004FFC0200364B2D800FFA";
    attribute INIT_39 of inst : label is "57904908011C248602386C0F284390AE092801648123C60A478C132019005D81";
    attribute INIT_3A of inst : label is "01007FFFE8080D9156AAA802101142812740A03A050280294800A14494002234";
    attribute INIT_3B of inst : label is "012001FFFD0150101F41087FFE00286100850000803EA248425FFF110408C108";
    attribute INIT_3C of inst : label is "B8BB5C59AE3AE6B8B35C59AE2CD7166B8B35C59AE2DB2496E014024001B24B6E";
    attribute INIT_3D of inst : label is "0A4201826400000002FFD40111803200E2AE2CD7176B8BB5C5D7173AE2ED7176";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000C8F1F74FC838";
    attribute INIT_3F of inst : label is "3E00000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "72492E492C92684B2B944B6185972896C3261C4F5E187048D603000000000121";
    attribute INIT_01 of inst : label is "EDFF38F088766114422699312484C836289D1249E49AE08E42C8C49124448952";
    attribute INIT_02 of inst : label is "9892CBDC8C2E464427842AED347D503EA9238F248248D9B05F91393263246985";
    attribute INIT_03 of inst : label is "198ED10A588D621892BC452114888891124C85B44B59389A218F68967C9C080C";
    attribute INIT_04 of inst : label is "3C849158C00AE2649274A4A5827EA0C269731533FFC166030833218840C0404C";
    attribute INIT_05 of inst : label is "9D0681925D2409249AC52428C6991E1DB3CF680AA7864D802200440281140082";
    attribute INIT_06 of inst : label is "0989831C36981809B7442182925509B4C4C84CCD86644A24499849A044492699";
    attribute INIT_07 of inst : label is "83330DB324E1B39AD8D289420942462504C89D5B6F093320693270C296111F18";
    attribute INIT_08 of inst : label is "E327A1039DD02B6619ADA5EC224263130E463D14114109140C21003434184049";
    attribute INIT_09 of inst : label is "418312322484924CA423389111A68A0921A7141360828C8919109249265C9004";
    attribute INIT_0A of inst : label is "911222492493341264CB666278D856159024981B109016D8080D326849061216";
    attribute INIT_0B of inst : label is "76108A92A4828C3082E03241C0448C99C49B842219219264EB9749DC710F3C91";
    attribute INIT_0C of inst : label is "210622011C111149013B21921928482486461192CC3A0C32118CB4310C8C25C2";
    attribute INIT_0D of inst : label is "19209A026982D20A4CDFF70080810F84209F2996574D21A4710184800C111148";
    attribute INIT_0E of inst : label is "8382180E41BC9264D9E2E4C8BA43610E73683C21BFE68F0864661C2949C6061C";
    attribute INIT_0F of inst : label is "B465A422229F26C9F26C311E40617B4C1133280E6200BDAF1AD3592D99063233";
    attribute INIT_10 of inst : label is "32480852202493924DA440492E241C48C7125B12306E241C48C7125B1230754C";
    attribute INIT_11 of inst : label is "9986186B06682344336135202D0D7090C609230E224C9E04C49391C258D02618";
    attribute INIT_12 of inst : label is "844FF30223000FF8880B6C5158374028DC566166071C9496849E269069C3594E";
    attribute INIT_13 of inst : label is "0592060449AE46709FDEED08E920007DDA02193264011F3C6849ED35EDD4CDF0";
    attribute INIT_14 of inst : label is "0A854B1493143BDE3A4603E1899B64A0F8E3E260DD06548B4924FE40743B3525";
    attribute INIT_15 of inst : label is "364C849E6EB4726846B0228202292664D660278126DFCC6B619827408DF9DE11";
    attribute INIT_16 of inst : label is "319B3C22D28690A673384C1819942B3BFCA121A60450484452493A4BC482D932";
    attribute INIT_17 of inst : label is "5149AA28A59000350031E0343C20CB0924D33843040E3000E64B59C174C13822";
    attribute INIT_18 of inst : label is "46664848166F1AC4D2CC4C4809BFF5A09719CC7318E6D831002C5632C65E3354";
    attribute INIT_19 of inst : label is "274CC784701249DB24D9E116942648E200080806B21884347649B499C886F3B2";
    attribute INIT_1A of inst : label is "80CDA6810BADC00241C3106260506643D238E38E3031F4C80888CCCC82232223";
    attribute INIT_1B of inst : label is "32424248C4904F16C486D192329B737C04C0000000000000000001F506F801B0";
    attribute INIT_1C of inst : label is "3318C4411C88448162773849388851D9E26DC70C0FF8E018600CE199040A4191";
    attribute INIT_1D of inst : label is "1CD8249CA4C527D9DB7463779B1022311A6E1992DECC93975939AF116CD6E627";
    attribute INIT_1E of inst : label is "F09210490C1F39242784091143689524E609064848CE480CC919066866036CD2";
    attribute INIT_1F of inst : label is "00100000100007F80007F8000000078000000000000000000000FFABAEBFBFAE";
    attribute INIT_20 of inst : label is "0707000300000000000000000000000000000000000000000000008004000008";
    attribute INIT_21 of inst : label is "00000002222AAAAAAAAAAA02022A8A8A8A8A8A8A828207070700070307070007";
    attribute INIT_22 of inst : label is "000000000000000000000000000001FFFFFF00FF8B8D75031000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "B6DB4D24920E4A3638D892E0A142E23F7E38B585B8D1B3DA991734ADC2B49B5E";
    attribute INIT_25 of inst : label is "09E6B163483F126123F9FC6C2D42C4AE238473188E1735BFEFF0C878EBFED24D";
    attribute INIT_26 of inst : label is "0B7E19FB605884828FDFCFE7F0B616A09E6A1621F7E59205A8FDFEFF7F8B716B";
    attribute INIT_27 of inst : label is "0182100180460C6EC077DFDCC0C0E2D6C90BBB7E111D3F6979030B0A3F1F7F0B";
    attribute INIT_28 of inst : label is "12082A80C200A80123C0020000CD1542155992499992499914924CC22AA28AA0";
    attribute INIT_29 of inst : label is "40A200AAA800140AAAAAAAAAAAAA803C991FE260000C04809080824273F83060";
    attribute INIT_2A of inst : label is "AA05555020445444445501111102AAAAAAAAAAAAAAAAAAAAAA81111111020444";
    attribute INIT_2B of inst : label is "5555502AAAAAAAAAAAA0AA80000000000000000000000000000004101040AAAA";
    attribute INIT_2C of inst : label is "000000000000000000FC15105440545411150150511114414102222222220555";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "000000000666477177066040442200111111111110000020202881191E4AC6A4";
    attribute INIT_31 of inst : label is "000000008E86E7D58EE0E242A0A8AA80888AAA268FFF7471F5FFBFF7F3FF5FD3";
    attribute INIT_32 of inst : label is "000000002E8EEE4E2C6A8A2AAAA8A6EF3344626040422EECE6EEE2EC6AE4CCC0";
    attribute INIT_33 of inst : label is "0000000004404444408888088088808A88ABB93B303B744EAAA822222A880880";
    attribute INIT_34 of inst : label is "000000005FFFFFFBFFCEEEEEEE228AB199DD9BB11115113BBBBBBBBBBFCFFFFF";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "4980F6E6761918B60E293149119246496496496496490FFF627476D92CE6DFF8";
    attribute INIT_39 of inst : label is "53B04871E0CC2439C198666A031B062C29160164092020124040262931484CCD";
    attribute INIT_3A of inst : label is "831000003888C111540000031680501092082490411389231891E3019C482214";
    attribute INIT_3B of inst : label is "A47208000711711181D3190004000C01083719098C83008CC400018046401198";
    attribute INIT_3C of inst : label is "AC93D649EB3EE3AC93D649EB24F5927AC93D649EB2492496CA4148E419B6D924";
    attribute INIT_3D of inst : label is "12822104C524000000001C6519852624B3EB24F5927AC93D67F5927EB24F5927";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000C808FDCDC824";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
