-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "105AE6667FF9AFF2676E2472C2C159240F03F4D949870000A63C36C5A7969A33";
    attribute INIT_01 of inst : label is "FFFFFF06DA849F0E49CA20C861FE4C677717FFFFB6D36D37D264A108797012FF";
    attribute INIT_02 of inst : label is "2CB0471220AC484116A2915498041008082011CF7DDAF3EF4C9933693F3BF577";
    attribute INIT_03 of inst : label is "A7FED0FEF34E1923F9265DF4283EC770B88EE91BAE32E29FF94C9B260390FFBB";
    attribute INIT_04 of inst : label is "7A5CF73CF3C18306601830660FD3CCC043643021EEEBE6DDCFFC7F7F4E3D7EF7";
    attribute INIT_05 of inst : label is "7FF9F634A64024921E4D48C26FEA037FFDFE73C3A7DFBF7E7677B76FFA6D6D3B";
    attribute INIT_06 of inst : label is "6561036B76B76B76B7A89E4E7C1FC0854AE03EE01FE037E01E34D3F7FC8653CA";
    attribute INIT_07 of inst : label is "FD7BB5FEBF84720E12B341505DB787BBC0A523F6992E4A497252D5859584B561";
    attribute INIT_08 of inst : label is "6842C128C5B50CD29FE1243FFEB5759C8F67A3C60BE2BE0BE2BAF99F4529EBC3";
    attribute INIT_09 of inst : label is "669A604499D99DAA068FB5290FDB0F3411DF836A6337584E201724014C9DDD0D";
    attribute INIT_0A of inst : label is "18C69268FB5272C6FFF5F504FBFEE7BC738CF36DFB7284370BCEFFFFAAAAFE9A";
    attribute INIT_0B of inst : label is "CD4F008276FB1DBCB9F5EB31EBB1EB31EBBEF7DF6C51CDE1998A0CB8F5D87FDC";
    attribute INIT_0C of inst : label is "392C6923E6F52557E88710F8EC74BA80F59312B414D723F044889626224AA922";
    attribute INIT_0D of inst : label is "23FFFFFFFFCC87FDD777EBBCD92C4493249D1BBF4CFE745D9092E865FF96FBF6";
    attribute INIT_0E of inst : label is "7A8013074C18FB34D2129E0E0B965C52A4DE7F965F7EF54FE6D62EECF80789FD";
    attribute INIT_0F of inst : label is "0001545555216AA912A82CC89A691E958EE4C81B41420AAD05082AAA46EDE62C";
    attribute INIT_10 of inst : label is "105AE6667FF9AFF2676E2472C2C159240F03F4D949870000A63C36C5A7969A33";
    attribute INIT_11 of inst : label is "FFFFFF06DA849F0E49CA20C861FE4C677717FFFFB6D36D37D264A108797012FF";
    attribute INIT_12 of inst : label is "2CB0471220AC484116A2915498041008082011CF7DDAF3EF4C9933693F3BF577";
    attribute INIT_13 of inst : label is "A7FED0FEF34E1923F9265DF4283EC770B88EE91BAE32E29FF94C9B260390FFBB";
    attribute INIT_14 of inst : label is "7A5CF73CF3C18306601830660FD3CCC043643021EEEBE6DDCFFC7F7F4E3D7EF7";
    attribute INIT_15 of inst : label is "7FF9F634A64024921E4D48C26FEA037FFDFE73C3A7DFBF7E7677B76FFA6D6D3B";
    attribute INIT_16 of inst : label is "6561036B76B76B76B7A89E4E7C1FC0854AE03EE01FE037E01E34D3F7FC8653CA";
    attribute INIT_17 of inst : label is "FD7BB5FEBF84720E12B341505DB787BBC0A523F6992E4A497252D5859584B561";
    attribute INIT_18 of inst : label is "6842C128C5B50CD29FE1243FFEB5759C8F67A3C60BE2BE0BE2BAF99F4529EBC3";
    attribute INIT_19 of inst : label is "669A604499D99DAA068FB5290FDB0F3411DF836A6337584E201724014C9DDD0D";
    attribute INIT_1A of inst : label is "18C69268FB5272C6FFF5F504FBFEE7BC738CF36DFB7284370BCEFFFFAAAAFE9A";
    attribute INIT_1B of inst : label is "CD4F008276FB1DBCB9F5EB31EBB1EB31EBBEF7DF6C51CDE1998A0CB8F5D87FDC";
    attribute INIT_1C of inst : label is "392C6923E6F52557E88710F8EC74BA80F59312B414D723F044889626224AA922";
    attribute INIT_1D of inst : label is "23FFFFFFFFCC87FDD777EBBCD92C4493249D1BBF4CFE745D9092E865FF96FBF6";
    attribute INIT_1E of inst : label is "7A8013074C18FB34D2129E0E0B965C52A4DE7F965F7EF54FE6D62EECF80789FD";
    attribute INIT_1F of inst : label is "0001545555216AA912A82CC89A691E958EE4C81B41420AAD05082AAA46EDE62C";
    attribute INIT_20 of inst : label is "D8FD82A00425F9D9CFFF84BB4773DF049347931CE20A3A84AE2090E309440410";
    attribute INIT_21 of inst : label is "83110001000100101380A0282544002C24242CD0F9C3F38752AA0AB6D5E994AF";
    attribute INIT_22 of inst : label is "7DD66BACD7EEB2ED7ACBB5E9349102C7C4D924B25000000000048A288D56053A";
    attribute INIT_23 of inst : label is "554EE7EA6FD9015173753B9DD4EE6753B9D365994F97F9C9FFD94A466D77F2D7";
    attribute INIT_24 of inst : label is "37BBC548C741FF6A9A83FFFFFF8FAE604E8A1108508B6C5441155146F8CC8601";
    attribute INIT_25 of inst : label is "490002010482402482231129AEB2B8EEF72B5DAE54EEF76623BBDC4546773BC1";
    attribute INIT_26 of inst : label is "7BF7AE5543BBDDD19DCEBAB4E81111112109889084C46E004124492480000000";
    attribute INIT_27 of inst : label is "FFFFFFFFF8E5012282AFD0B0BF4022908A4011C0C43E1933505040CA08220118";
    attribute INIT_28 of inst : label is "D8FD82A00425F9D9CFFF84BB4773DF049347931CE20A3A84AE2090E309440410";
    attribute INIT_29 of inst : label is "83110001000100101380A0282544002C24242CD0F9C3F38752AA0AB6D5E994AF";
    attribute INIT_2A of inst : label is "7DD66BACD7EEB2ED7ACBB5E9349102C7C4D924B25000000000048A288D56053A";
    attribute INIT_2B of inst : label is "554EE7EA6FD9015173753B9DD4EE6753B9D365994F97F9C9FFD94A466D77F2D7";
    attribute INIT_2C of inst : label is "37BBC548C741FF6A9A83FFFFFF8FAE604E8A1108508B6C5441155146F8CC8601";
    attribute INIT_2D of inst : label is "490002010482402482231129AEB2B8EEF72B5DAE54EEF76623BBDC4546773BC1";
    attribute INIT_2E of inst : label is "7BF7AE5543BBDDD19DCEBAB4E81111112109889084C46E004124492480000000";
    attribute INIT_2F of inst : label is "FFFFFFFFF8E5012282AFD0B0BF4022908A4011C0C43E1933505040CA08220118";
    attribute INIT_30 of inst : label is "D8FD82A00425F9D9CFFF84BB4773DF049347931CE20A3A84AE2090E309440410";
    attribute INIT_31 of inst : label is "83110001000100101380A0282544002C24242CD0F9C3F38752AA0AB6D5E994AF";
    attribute INIT_32 of inst : label is "7DD66BACD7EEB2ED7ACBB5E9349102C7C4D924B25000000000048A288D56053A";
    attribute INIT_33 of inst : label is "554EE7EA6FD9015173753B9DD4EE6753B9D365994F97F9C9FFD94A466D77F2D7";
    attribute INIT_34 of inst : label is "37BBC548C741FF6A9A83FFFFFF8FAE604E8A1108508B6C5441155146F8CC8601";
    attribute INIT_35 of inst : label is "490002010482402482231129AEB2B8EEF72B5DAE54EEF76623BBDC4546773BC1";
    attribute INIT_36 of inst : label is "7BF7AE5543BBDDD19DCEBAB4E81111112109889084C46E004124492480000000";
    attribute INIT_37 of inst : label is "FFFFFFFFF8E5012282AFD0B0BF4022908A4011C0C43E1933505040CA08220118";
    attribute INIT_38 of inst : label is "D8FD82A00425F9D9CFFF84BB4773DF049347931CE20A3A84AE2090E309440410";
    attribute INIT_39 of inst : label is "83110001000100101380A0282544002C24242CD0F9C3F38752AA0AB6D5E994AF";
    attribute INIT_3A of inst : label is "7DD66BACD7EEB2ED7ACBB5E9349102C7C4D924B25000000000048A288D56053A";
    attribute INIT_3B of inst : label is "554EE7EA6FD9015173753B9DD4EE6753B9D365994F97F9C9FFD94A466D77F2D7";
    attribute INIT_3C of inst : label is "37BBC548C741FF6A9A83FFFFFF8FAE604E8A1108508B6C5441155146F8CC8601";
    attribute INIT_3D of inst : label is "490002010482402482231129AEB2B8EEF72B5DAE54EEF76623BBDC4546773BC1";
    attribute INIT_3E of inst : label is "7BF7AE5543BBDDD19DCEBAB4E81111112109889084C46E004124492480000000";
    attribute INIT_3F of inst : label is "FFFFFFFFF8E5012282AFD0B0BF4022908A4011C0C43E1933505040CA08220118";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "EBA000000040D40D5FB9D9F4C4C9814B2806000083C80000CC5A95639433A36A";
    attribute INIT_01 of inst : label is "FFFFFE010E9B90A370DB6C270C81AB59DD83FC24CA28820A299BDBD6FA2D0494";
    attribute INIT_02 of inst : label is "451AF9834700CE8A2A2DC28BCE298324530649F0D2FD9197A922AF38142D0A4F";
    attribute INIT_03 of inst : label is "4FFC9D4332400661B21163DBD229DA88A5B71BFE4BA4B9200099709158647F01";
    attribute INIT_04 of inst : label is "588140F14F0B3264C4B3264C68A06BBB719DBBFA06952F41511200D8A98480C8";
    attribute INIT_05 of inst : label is "031212C848B64B2C8D01AD2D84DB6CA822510610E41000400008491448236C0B";
    attribute INIT_06 of inst : label is "8282688C48C48C48C45F4EA83EAFAEE99289A689A789878982599716CA3139A7";
    attribute INIT_07 of inst : label is "91E482C8F04999B19184CA22121828240C4990D9269184B488251A1A0A094686";
    attribute INIT_08 of inst : label is "672B166B12F4816A510E55A6FCDCC82B54AA4568960B60B60963F0B04C12CD0D";
    attribute INIT_09 of inst : label is "084B0919110B307F0036D252003840A181216641426DFF83C72452C1C40C6425";
    attribute INIT_0A of inst : label is "AF68490301243FF3FFEA0440BAE2288E3CA1D9EF751D07D140A155550000F84B";
    attribute INIT_0B of inst : label is "C40766D09186327AA416925EB25E92DEB2C96CFBFE1E60A43666C16F09000796";
    attribute INIT_0C of inst : label is "104195D44903C3DACC5CA385B5C90B40E400A7F603240C4E187705C14F87700F";
    attribute INIT_0D of inst : label is "2FFFFFFFFF1257F81A493AD3D648E8680327EAF883FC9F962566170CFF401E0B";
    attribute INIT_0E of inst : label is "1C00066D19B3606E356D216196A289BF3B6530A28A51C1E3CB2974A8C323C662";
    attribute INIT_0F of inst : label is "0001CC333CA0C658919C18010487812DF48B73222D4B2AC8B56CA935B902C153";
    attribute INIT_10 of inst : label is "EBA000000040D40D5FB9D9F4C4C9814B2806000083C80000CC5A95639433A36A";
    attribute INIT_11 of inst : label is "FFFFFE010E9B90A370DB6C270C81AB59DD83FC24CA28820A299BDBD6FA2D0494";
    attribute INIT_12 of inst : label is "451AF9834700CE8A2A2DC28BCE298324530649F0D2FD9197A922AF38142D0A4F";
    attribute INIT_13 of inst : label is "4FFC9D4332400661B21163DBD229DA88A5B71BFE4BA4B9200099709158647F01";
    attribute INIT_14 of inst : label is "588140F14F0B3264C4B3264C68A06BBB719DBBFA06952F41511200D8A98480C8";
    attribute INIT_15 of inst : label is "031212C848B64B2C8D01AD2D84DB6CA822510610E41000400008491448236C0B";
    attribute INIT_16 of inst : label is "8282688C48C48C48C45F4EA83EAFAEE99289A689A789878982599716CA3139A7";
    attribute INIT_17 of inst : label is "91E482C8F04999B19184CA22121828240C4990D9269184B488251A1A0A094686";
    attribute INIT_18 of inst : label is "672B166B12F4816A510E55A6FCDCC82B54AA4568960B60B60963F0B04C12CD0D";
    attribute INIT_19 of inst : label is "084B0919110B307F0036D252003840A181216641426DFF83C72452C1C40C6425";
    attribute INIT_1A of inst : label is "AF68490301243FF3FFEA0440BAE2288E3CA1D9EF751D07D140A155550000F84B";
    attribute INIT_1B of inst : label is "C40766D09186327AA416925EB25E92DEB2C96CFBFE1E60A43666C16F09000796";
    attribute INIT_1C of inst : label is "104195D44903C3DACC5CA385B5C90B40E400A7F603240C4E187705C14F87700F";
    attribute INIT_1D of inst : label is "2FFFFFFFFF1257F81A493AD3D648E8680327EAF883FC9F962566170CFF401E0B";
    attribute INIT_1E of inst : label is "1C00066D19B3606E356D216196A289BF3B6530A28A51C1E3CB2974A8C323C662";
    attribute INIT_1F of inst : label is "0001CC333CA0C658919C18010487812DF48B73222D4B2AC8B56CA935B902C153";
    attribute INIT_20 of inst : label is "19B1917CD351029290069929AA802CCB394B1A539D9A4FBB59C95A9A448B335D";
    attribute INIT_21 of inst : label is "112323222322233320F3DE8D00DC200C000008D822184433CBC56249601ADABB";
    attribute INIT_22 of inst : label is "8B2C86DB241965B205B649124964F7FC211B24967288C8C8C8CC012400036FBF";
    attribute INIT_23 of inst : label is "58E098055866D697A58A423A2900E9A423E44DE28333FA19FF9D75ACED261C8C";
    attribute INIT_24 of inst : label is "544234BBBC5AFF76CDBAFFFFFF181A85D2B1A66B4B314148F7676C610456CC98";
    attribute INIT_25 of inst : label is "0820100800100804007868C64A2E2D7118AC92896D5108E855C46348AA884480";
    attribute INIT_26 of inst : label is "860C6948B584422AE231244C9E0303030001818000C0F2004820010410410082";
    attribute INIT_27 of inst : label is "FFFFFFFFFF4FF134708D5460351B3BBBB6EC83120D1F8851367380EE502B281A";
    attribute INIT_28 of inst : label is "19B1917CD351029290069929AA802CCB394B1A539D9A4FBB59C95A9A448B335D";
    attribute INIT_29 of inst : label is "112323222322233320F3DE8D00DC200C000008D822184433CBC56249601ADABB";
    attribute INIT_2A of inst : label is "8B2C86DB241965B205B649124964F7FC211B24967288C8C8C8CC012400036FBF";
    attribute INIT_2B of inst : label is "58E098055866D697A58A423A2900E9A423E44DE28333FA19FF9D75ACED261C8C";
    attribute INIT_2C of inst : label is "544234BBBC5AFF76CDBAFFFFFF181A85D2B1A66B4B314148F7676C610456CC98";
    attribute INIT_2D of inst : label is "0820100800100804007868C64A2E2D7118AC92896D5108E855C46348AA884480";
    attribute INIT_2E of inst : label is "860C6948B584422AE231244C9E0303030001818000C0F2004820010410410082";
    attribute INIT_2F of inst : label is "FFFFFFFFFF4FF134708D5460351B3BBBB6EC83120D1F8851367380EE502B281A";
    attribute INIT_30 of inst : label is "19B1917CD351029290069929AA802CCB394B1A539D9A4FBB59C95A9A448B335D";
    attribute INIT_31 of inst : label is "112323222322233320F3DE8D00DC200C000008D822184433CBC56249601ADABB";
    attribute INIT_32 of inst : label is "8B2C86DB241965B205B649124964F7FC211B24967288C8C8C8CC012400036FBF";
    attribute INIT_33 of inst : label is "58E098055866D697A58A423A2900E9A423E44DE28333FA19FF9D75ACED261C8C";
    attribute INIT_34 of inst : label is "544234BBBC5AFF76CDBAFFFFFF181A85D2B1A66B4B314148F7676C610456CC98";
    attribute INIT_35 of inst : label is "0820100800100804007868C64A2E2D7118AC92896D5108E855C46348AA884480";
    attribute INIT_36 of inst : label is "860C6948B584422AE231244C9E0303030001818000C0F2004820010410410082";
    attribute INIT_37 of inst : label is "FFFFFFFFFF4FF134708D5460351B3BBBB6EC83120D1F8851367380EE502B281A";
    attribute INIT_38 of inst : label is "19B1917CD351029290069929AA802CCB394B1A539D9A4FBB59C95A9A448B335D";
    attribute INIT_39 of inst : label is "112323222322233320F3DE8D00DC200C000008D822184433CBC56249601ADABB";
    attribute INIT_3A of inst : label is "8B2C86DB241965B205B649124964F7FC211B24967288C8C8C8CC012400036FBF";
    attribute INIT_3B of inst : label is "58E098055866D697A58A423A2900E9A423E44DE28333FA19FF9D75ACED261C8C";
    attribute INIT_3C of inst : label is "544234BBBC5AFF76CDBAFFFFFF181A85D2B1A66B4B314148F7676C610456CC98";
    attribute INIT_3D of inst : label is "0820100800100804007868C64A2E2D7118AC92896D5108E855C46348AA884480";
    attribute INIT_3E of inst : label is "860C6948B584422AE231244C9E0303030001818000C0F2004820010410410082";
    attribute INIT_3F of inst : label is "FFFFFFFFFF4FF134708D5460351B3BBBB6EC83120D1F8851367380EE502B281A";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "00908CCCF078537977D5EE862E0CC8466C03054083C7AAAA1181481848484484";
    attribute INIT_01 of inst : label is "FFFFFE38000738FE78DB72338E6F2E611107FCF5C5145142A064C3E0FB6E0679";
    attribute INIT_02 of inst : label is "F59CFA53813446020AA134936812689A24D1350255DBB0BA8C58BA3845B97277";
    attribute INIT_03 of inst : label is "77FD4CE2EEC60D80733439331C14A720514C45C336BB69C948EBF5BD9ED87F73";
    attribute INIT_04 of inst : label is "B5AC4BA61034C9D3BB4C9D3BA0A9E66361341A1801532F8EDD133A5E2C886432";
    attribute INIT_05 of inst : label is "96CEA64E734026D20D692E2A4FDB447B45ADB0612952A50A1D1631D47033B60D";
    attribute INIT_06 of inst : label is "B2F30A4824864824864C13B845EFB26165D185D180D180D18036B431DDB8ED9D";
    attribute INIT_07 of inst : label is "F5F9B2FAFE8EA61C94648A761E9D6AB9647000F7C5F5672FAF39CACACBCC72B2";
    attribute INIT_08 of inst : label is "4948652A65A506CA8CB31519FCA0F11C8E47B3DA26A06A06A06B5089451CE5E5";
    attribute INIT_09 of inst : label is "2082214E6C96C9550097B3BC05DF85A511D6A24A63A963A266279241AC2C75AD";
    attribute INIT_0A of inst : label is "A10A924973395E41FFEAAEEFAAA0A82E28E9DDC4505C050540EB50505050F882";
    attribute INIT_0B of inst : label is "C508C6B115FA3DB639F9C3A9C3A9E3A9E3A77A41259040CADCC6464B59E87F80";
    attribute INIT_0C of inst : label is "175C65CF9957235CC04AB16EADBA8B00E50EF5560750BD89D4440B1DEE4660EE";
    attribute INIT_0D of inst : label is "A3FFFFFFFF6CDBFADC72EBAEDC643EEAB779E338A7FDE798D1DA4926FF6BD7A6";
    attribute INIT_0E of inst : label is "9E000993E64C57AAAF29C3AB06FAC82104AF7DFACDEDC597DFCAEE12F003C726";
    attribute INIT_0F of inst : label is "0001FC0F0C03E1C5947D168377D6D6884E6CA4C325516A0C9505A8518F8FDDE3";
    attribute INIT_10 of inst : label is "00908CCCF078537977D5EE862E0CC8466C03054083C7AAAA1181481848484484";
    attribute INIT_11 of inst : label is "FFFFFE38000738FE78DB72338E6F2E611107FCF5C5145142A064C3E0FB6E0679";
    attribute INIT_12 of inst : label is "F59CFA53813446020AA134936812689A24D1350255DBB0BA8C58BA3845B97277";
    attribute INIT_13 of inst : label is "77FD4CE2EEC60D80733439331C14A720514C45C336BB69C948EBF5BD9ED87F73";
    attribute INIT_14 of inst : label is "B5AC4BA61034C9D3BB4C9D3BA0A9E66361341A1801532F8EDD133A5E2C886432";
    attribute INIT_15 of inst : label is "96CEA64E734026D20D692E2A4FDB447B45ADB0612952A50A1D1631D47033B60D";
    attribute INIT_16 of inst : label is "B2F30A4824864824864C13B845EFB26165D185D180D180D18036B431DDB8ED9D";
    attribute INIT_17 of inst : label is "F5F9B2FAFE8EA61C94648A761E9D6AB9647000F7C5F5672FAF39CACACBCC72B2";
    attribute INIT_18 of inst : label is "4948652A65A506CA8CB31519FCA0F11C8E47B3DA26A06A06A06B5089451CE5E5";
    attribute INIT_19 of inst : label is "2082214E6C96C9550097B3BC05DF85A511D6A24A63A963A266279241AC2C75AD";
    attribute INIT_1A of inst : label is "A10A924973395E41FFEAAEEFAAA0A82E28E9DDC4505C050540EB50505050F882";
    attribute INIT_1B of inst : label is "C508C6B115FA3DB639F9C3A9C3A9E3A9E3A77A41259040CADCC6464B59E87F80";
    attribute INIT_1C of inst : label is "175C65CF9957235CC04AB16EADBA8B00E50EF5560750BD89D4440B1DEE4660EE";
    attribute INIT_1D of inst : label is "A3FFFFFFFF6CDBFADC72EBAEDC643EEAB779E338A7FDE798D1DA4926FF6BD7A6";
    attribute INIT_1E of inst : label is "9E000993E64C57AAAF29C3AB06FAC82104AF7DFACDEDC597DFCAEE12F003C726";
    attribute INIT_1F of inst : label is "0001FC0F0C03E1C5947D168377D6D6884E6CA4C325516A0C9505A8518F8FDDE3";
    attribute INIT_20 of inst : label is "D0890930E306294B5AFE9923BE993B16D650CB9D5EAA810857EA5CE38403238C";
    attribute INIT_21 of inst : label is "E75555444455555557C5C41C48FC444C484848FC195C32FA930972A495CB0288";
    attribute INIT_22 of inst : label is "95E7BB4D5EED34F5EEF3D7AFD7AC9871231B659644555511551110451543BC5C";
    attribute INIT_23 of inst : label is "416A76C9515914D5087368BFCDA2FE36ABB20DB8D933FB59FF9B7338DF24E5C7";
    attribute INIT_24 of inst : label is "3D0E9448A047FF421082FFFFFF2924284481888A44444440230167039058151A";
    attribute INIT_25 of inst : label is "D36936936DA6D36DB6804DCEC38FCCD42A2844F14CE432741310894026211040";
    attribute INIT_26 of inst : label is "1A3B0C4033D0E8C988443834EE0E0E0E18C6070C630382249B491269B49A4926";
    attribute INIT_27 of inst : label is "FFFFFFFFFD98047340A575DD6F227F9C06F240D1C51FC8132151CDEA336A18BA";
    attribute INIT_28 of inst : label is "D0890930E306294B5AFE9923BE993B16D650CB9D5EAA810857EA5CE38403238C";
    attribute INIT_29 of inst : label is "E75555444455555557C5C41C48FC444C484848FC195C32FA930972A495CB0288";
    attribute INIT_2A of inst : label is "95E7BB4D5EED34F5EEF3D7AFD7AC9871231B659644555511551110451543BC5C";
    attribute INIT_2B of inst : label is "416A76C9515914D5087368BFCDA2FE36ABB20DB8D933FB59FF9B7338DF24E5C7";
    attribute INIT_2C of inst : label is "3D0E9448A047FF421082FFFFFF2924284481888A44444440230167039058151A";
    attribute INIT_2D of inst : label is "D36936936DA6D36DB6804DCEC38FCCD42A2844F14CE432741310894026211040";
    attribute INIT_2E of inst : label is "1A3B0C4033D0E8C988443834EE0E0E0E18C6070C630382249B491269B49A4926";
    attribute INIT_2F of inst : label is "FFFFFFFFFD98047340A575DD6F227F9C06F240D1C51FC8132151CDEA336A18BA";
    attribute INIT_30 of inst : label is "D0890930E306294B5AFE9923BE993B16D650CB9D5EAA810857EA5CE38403238C";
    attribute INIT_31 of inst : label is "E75555444455555557C5C41C48FC444C484848FC195C32FA930972A495CB0288";
    attribute INIT_32 of inst : label is "95E7BB4D5EED34F5EEF3D7AFD7AC9871231B659644555511551110451543BC5C";
    attribute INIT_33 of inst : label is "416A76C9515914D5087368BFCDA2FE36ABB20DB8D933FB59FF9B7338DF24E5C7";
    attribute INIT_34 of inst : label is "3D0E9448A047FF421082FFFFFF2924284481888A44444440230167039058151A";
    attribute INIT_35 of inst : label is "D36936936DA6D36DB6804DCEC38FCCD42A2844F14CE432741310894026211040";
    attribute INIT_36 of inst : label is "1A3B0C4033D0E8C988443834EE0E0E0E18C6070C630382249B491269B49A4926";
    attribute INIT_37 of inst : label is "FFFFFFFFFD98047340A575DD6F227F9C06F240D1C51FC8132151CDEA336A18BA";
    attribute INIT_38 of inst : label is "D0890930E306294B5AFE9923BE993B16D650CB9D5EAA810857EA5CE38403238C";
    attribute INIT_39 of inst : label is "E75555444455555557C5C41C48FC444C484848FC195C32FA930972A495CB0288";
    attribute INIT_3A of inst : label is "95E7BB4D5EED34F5EEF3D7AFD7AC9871231B659644555511551110451543BC5C";
    attribute INIT_3B of inst : label is "416A76C9515914D5087368BFCDA2FE36ABB20DB8D933FB59FF9B7338DF24E5C7";
    attribute INIT_3C of inst : label is "3D0E9448A047FF421082FFFFFF2924284481888A44444440230167039058151A";
    attribute INIT_3D of inst : label is "D36936936DA6D36DB6804DCEC38FCCD42A2844F14CE432741310894026211040";
    attribute INIT_3E of inst : label is "1A3B0C4033D0E8C988443834EE0E0E0E18C6070C630382249B491269B49A4926";
    attribute INIT_3F of inst : label is "FFFFFFFFFD98047340A575DD6F227F9C06F240D1C51FC8132151CDEA336A18BA";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "F190AEEED4401B712F9DEC85070BCC6EEE028448C188CCCC0000000000000000";
    attribute INIT_01 of inst : label is "FFFFFFB888824070550D3E61A66E253CAA83FE776410410BA240C17078D716EF";
    attribute INIT_02 of inst : label is "A49C93D1E13456C30E8EB0C3EA492248924491067B016018E7DC9E280F1FF33F";
    attribute INIT_03 of inst : label is "6FFF4DB0CD801D90F98F1E231A06A5A85B4856A1F75F75BDEEDF9DBF1FD87F93";
    attribute INIT_04 of inst : label is "80DC17241066FD9F766FD9F77430345BF125129B0AD26281C20A0676259BF77B";
    attribute INIT_05 of inst : label is "BCF9F4746E4024930FCD26C3CF453050EB2C7841A2448912260D2B5E40029304";
    attribute INIT_06 of inst : label is "63234352F10B52B10F7DC073024FF26D556585E5856581E58026902BF59ADDDF";
    attribute INIT_07 of inst : label is "649923324C8FE60F0FF201FE1CB44FDFD76C0125C92ED6C976B6CC8C8D8D9363";
    attribute INIT_08 of inst : label is "D5ABC1B1C1388C8C2DE3985BFEB2BE556B955AA685E85E85E85950AD099B26C6";
    attribute INIT_09 of inst : label is "2FE1284DEED4CD910699235C0FD74F14D0FD8BA9A1F3BDC6579F1B70AC0CDF0A";
    attribute INIT_0A of inst : label is "15AEDB49B2360572FFD55050C20A5290B281FD6005210652828341414141FFE1";
    attribute INIT_0B of inst : label is "C140854134FB8F3651D959D559D559D559FCFB412590580BDDC5459D5DE82FCA";
    attribute INIT_0C of inst : label is "1D1C44FACCE622EEE85ED1EEFDEF8DC0F58AF65A1675A8DD547E8FF5EC45C8AD";
    attribute INIT_0D of inst : label is "0FFFFFFFFFC46BFFAE2EEDEEAF6C36CB365E4DFC40FF792FD9D24DA0FFCBFB34";
    attribute INIT_0E of inst : label is "AF0019DF677DB72286A5B7EE87D24C359793FDD24D2CE4B7FC4AEE21280385CE";
    attribute INIT_0F of inst : label is "0001FC00FBA3FFC00FF83EC055D29ECEABCD5D4FB68DB47EDA36D1D9F6CBF5E3";
    attribute INIT_10 of inst : label is "F190AEEED4401B712F9DEC85070BCC6EEE028448C188CCCC0000000000000000";
    attribute INIT_11 of inst : label is "FFFFFFB888824070550D3E61A66E253CAA83FE776410410BA240C17078D716EF";
    attribute INIT_12 of inst : label is "A49C93D1E13456C30E8EB0C3EA492248924491067B016018E7DC9E280F1FF33F";
    attribute INIT_13 of inst : label is "6FFF4DB0CD801D90F98F1E231A06A5A85B4856A1F75F75BDEEDF9DBF1FD87F93";
    attribute INIT_14 of inst : label is "80DC17241066FD9F766FD9F77430345BF125129B0AD26281C20A0676259BF77B";
    attribute INIT_15 of inst : label is "BCF9F4746E4024930FCD26C3CF453050EB2C7841A2448912260D2B5E40029304";
    attribute INIT_16 of inst : label is "63234352F10B52B10F7DC073024FF26D556585E5856581E58026902BF59ADDDF";
    attribute INIT_17 of inst : label is "649923324C8FE60F0FF201FE1CB44FDFD76C0125C92ED6C976B6CC8C8D8D9363";
    attribute INIT_18 of inst : label is "D5ABC1B1C1388C8C2DE3985BFEB2BE556B955AA685E85E85E85950AD099B26C6";
    attribute INIT_19 of inst : label is "2FE1284DEED4CD910699235C0FD74F14D0FD8BA9A1F3BDC6579F1B70AC0CDF0A";
    attribute INIT_1A of inst : label is "15AEDB49B2360572FFD55050C20A5290B281FD6005210652828341414141FFE1";
    attribute INIT_1B of inst : label is "C140854134FB8F3651D959D559D559D559FCFB412590580BDDC5459D5DE82FCA";
    attribute INIT_1C of inst : label is "1D1C44FACCE622EEE85ED1EEFDEF8DC0F58AF65A1675A8DD547E8FF5EC45C8AD";
    attribute INIT_1D of inst : label is "0FFFFFFFFFC46BFFAE2EEDEEAF6C36CB365E4DFC40FF792FD9D24DA0FFCBFB34";
    attribute INIT_1E of inst : label is "AF0019DF677DB72286A5B7EE87D24C359793FDD24D2CE4B7FC4AEE21280385CE";
    attribute INIT_1F of inst : label is "0001FC00FBA3FFC00FF83EC055D29ECEABCD5D4FB68DB47EDA36D1D9F6CBF5E3";
    attribute INIT_20 of inst : label is "A9DA9DF4DB7229495FADDCACA499B784960C8D4BDEACE5697DEA6E5950C23F4D";
    attribute INIT_21 of inst : label is "54454445454545454555541548F40440484848E49BED3F9A9D613077DCF3D23D";
    attribute INIT_22 of inst : label is "64925924B324926B7669ACDFAF94913D810B2C9266DDDDDD999DDE459FFD5595";
    attribute INIT_23 of inst : label is "9D6F66C901D014C747E17C93C5F24F17E93F8438ED1083C83FDFF628FB268592";
    attribute INIT_24 of inst : label is "21E8E1F3F09DFFD86639FFFFFF8BE560651DBCE19CE0859C2271BF41381E965A";
    attribute INIT_25 of inst : label is "000480492492492492410D8CCAAEA497ABC650A90897ABF6921E8F1D253D9E41";
    attribute INIT_26 of inst : label is "33BFE78C225EAF896F7796275800000000000000000002920000000002492490";
    attribute INIT_27 of inst : label is "FFFFFFFFF85FF08487D8A2A28822662D867240C0C41F4E1311134562014800AC";
    attribute INIT_28 of inst : label is "A9DA9DF4DB7229495FADDCACA499B784960C8D4BDEACE5697DEA6E5950C23F4D";
    attribute INIT_29 of inst : label is "54454445454545454555541548F40440484848E49BED3F9A9D613077DCF3D23D";
    attribute INIT_2A of inst : label is "64925924B324926B7669ACDFAF94913D810B2C9266DDDDDD999DDE459FFD5595";
    attribute INIT_2B of inst : label is "9D6F66C901D014C747E17C93C5F24F17E93F8438ED1083C83FDFF628FB268592";
    attribute INIT_2C of inst : label is "21E8E1F3F09DFFD86639FFFFFF8BE560651DBCE19CE0859C2271BF41381E965A";
    attribute INIT_2D of inst : label is "000480492492492492410D8CCAAEA497ABC650A90897ABF6921E8F1D253D9E41";
    attribute INIT_2E of inst : label is "33BFE78C225EAF896F7796275800000000000000000002920000000002492490";
    attribute INIT_2F of inst : label is "FFFFFFFFF85FF08487D8A2A28822662D867240C0C41F4E1311134562014800AC";
    attribute INIT_30 of inst : label is "A9DA9DF4DB7229495FADDCACA499B784960C8D4BDEACE5697DEA6E5950C23F4D";
    attribute INIT_31 of inst : label is "54454445454545454555541548F40440484848E49BED3F9A9D613077DCF3D23D";
    attribute INIT_32 of inst : label is "64925924B324926B7669ACDFAF94913D810B2C9266DDDDDD999DDE459FFD5595";
    attribute INIT_33 of inst : label is "9D6F66C901D014C747E17C93C5F24F17E93F8438ED1083C83FDFF628FB268592";
    attribute INIT_34 of inst : label is "21E8E1F3F09DFFD86639FFFFFF8BE560651DBCE19CE0859C2271BF41381E965A";
    attribute INIT_35 of inst : label is "000480492492492492410D8CCAAEA497ABC650A90897ABF6921E8F1D253D9E41";
    attribute INIT_36 of inst : label is "33BFE78C225EAF896F7796275800000000000000000002920000000002492490";
    attribute INIT_37 of inst : label is "FFFFFFFFF85FF08487D8A2A28822662D867240C0C41F4E1311134562014800AC";
    attribute INIT_38 of inst : label is "A9DA9DF4DB7229495FADDCACA499B784960C8D4BDEACE5697DEA6E5950C23F4D";
    attribute INIT_39 of inst : label is "54454445454545454555541548F40440484848E49BED3F9A9D613077DCF3D23D";
    attribute INIT_3A of inst : label is "64925924B324926B7669ACDFAF94913D810B2C9266DDDDDD999DDE459FFD5595";
    attribute INIT_3B of inst : label is "9D6F66C901D014C747E17C93C5F24F17E93F8438ED1083C83FDFF628FB268592";
    attribute INIT_3C of inst : label is "21E8E1F3F09DFFD86639FFFFFF8BE560651DBCE19CE0859C2271BF41381E965A";
    attribute INIT_3D of inst : label is "000480492492492492410D8CCAAEA497ABC650A90897ABF6921E8F1D253D9E41";
    attribute INIT_3E of inst : label is "33BFE78C225EAF896F7796275800000000000000000002920000000002492490";
    attribute INIT_3F of inst : label is "FFFFFFFFF85FF08487D8A2A28822662D867240C0C41F4E1311134562014800AC";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "E7A48222011110450F53D98D0D1C8AE661155818C32DF0F00000000000000000";
    attribute INIT_01 of inst : label is "FFFFFE40A15020225B0185029A08A1193313FC02C82082097C9B5C3704130090";
    attribute INIT_02 of inst : label is "0006C988D50AA4AAA8152EBA29924C93249926A9906DF2B02142842006040A0F";
    attribute INIT_03 of inst : label is "4FFCA9476FCC0480B2CB950B120308D00D10A060E10611250899504054487F20";
    attribute INIT_04 of inst : label is "95B0CC2080122648C800200438A0580370C21212980CC29405BE6991A3628442";
    attribute INIT_05 of inst : label is "92308848482D80000C93A30490810285A040C300DC912244824048920053B72D";
    attribute INIT_06 of inst : label is "4202C4E70E74A54A54134221260F9B4B9993ED93ED13E913E9C90D22C968A594";
    attribute INIT_07 of inst : label is "94A5124A52CB9D8A0004886700880A0D044A400A004104820C248909090B0242";
    attribute INIT_08 of inst : label is "9BD81A451A428129430A5286FDD89A2211289440D40D40D40D4114252A124404";
    attribute INIT_09 of inst : label is "08208C8901001005001042600468440280311405406163CACE205260A2010010";
    attribute INIT_0A of inst : label is "9398048120253DA4FFD55500A8A2609C8041C115513000138A4355005500F800";
    attribute INIT_0B of inst : label is "C124CC4E080C06400402204A204A204A2058201801863C2A6444410B5C082FE8";
    attribute INIT_0C of inst : label is "120A94B15411450AD039AA03138800C0E09CED4209A0554598A29499DA8A29CA";
    attribute INIT_0D of inst : label is "17FFFFFFFF146BF84A0930D3060AA028410720F8C9FC1C86254A2080FF048800";
    attribute INIT_0E of inst : label is "1400064C08100049242924E1D60002A1890410000240C06BCA6BE774D6C02026";
    attribute INIT_0F of inst : label is "00013C000FA3C04000040048E796212C50BA22A0262931409AA4C5042012D9CB";
    attribute INIT_10 of inst : label is "E7A48222011110450F53D98D0D1C8AE661155818C32DF0F00000000000000000";
    attribute INIT_11 of inst : label is "FFFFFE40A15020225B0185029A08A1193313FC02C82082097C9B5C3704130090";
    attribute INIT_12 of inst : label is "0006C988D50AA4AAA8152EBA29924C93249926A9906DF2B02142842006040A0F";
    attribute INIT_13 of inst : label is "4FFCA9476FCC0480B2CB950B120308D00D10A060E10611250899504054487F20";
    attribute INIT_14 of inst : label is "95B0CC2080122648C800200438A0580370C21212980CC29405BE6991A3628442";
    attribute INIT_15 of inst : label is "92308848482D80000C93A30490810285A040C300DC912244824048920053B72D";
    attribute INIT_16 of inst : label is "4202C4E70E74A54A54134221260F9B4B9993ED93ED13E913E9C90D22C968A594";
    attribute INIT_17 of inst : label is "94A5124A52CB9D8A0004886700880A0D044A400A004104820C248909090B0242";
    attribute INIT_18 of inst : label is "9BD81A451A428129430A5286FDD89A2211289440D40D40D40D4114252A124404";
    attribute INIT_19 of inst : label is "08208C8901001005001042600468440280311405406163CACE205260A2010010";
    attribute INIT_1A of inst : label is "9398048120253DA4FFD55500A8A2609C8041C115513000138A4355005500F800";
    attribute INIT_1B of inst : label is "C124CC4E080C06400402204A204A204A2058201801863C2A6444410B5C082FE8";
    attribute INIT_1C of inst : label is "120A94B15411450AD039AA03138800C0E09CED4209A0554598A29499DA8A29CA";
    attribute INIT_1D of inst : label is "17FFFFFFFF146BF84A0930D3060AA028410720F8C9FC1C86254A2080FF048800";
    attribute INIT_1E of inst : label is "1400064C08100049242924E1D60002A1890410000240C06BCA6BE774D6C02026";
    attribute INIT_1F of inst : label is "00013C000FA3C04000040048E796212C50BA22A0262931409AA4C5042012D9CB";
    attribute INIT_20 of inst : label is "1594504F92402B5B5FADBDC0809120F9203928433DF1C14851DF461862AA2249";
    attribute INIT_21 of inst : label is "40100001100110011111100103351808000101B04094812AA8DD51C2082A3A79";
    attribute INIT_22 of inst : label is "0945028A040A2880048201020108250832020900004000000000050800144201";
    attribute INIT_23 of inst : label is "3A9197D51226DA8B08113AB344E2CD138B350C36D63003D83F926DB092000B05";
    attribute INIT_24 of inst : label is "4A9552859028FFD96651FFFFFF561896925922252900012AA2AA0A828051E93C";
    attribute INIT_25 of inst : label is "924924924924924924AAA853C12D2D1A4D14904BAD1A4D695429152AA952A800";
    attribute INIT_26 of inst : label is "0444812AA429142A74BA85481B656565CE72B2E7395957249249924924924924";
    attribute INIT_27 of inst : label is "FFFFFFFFFA88200A0A0A0A00A0003328D4600A0A288100847BA3B4B54D2DA0D1";
    attribute INIT_28 of inst : label is "1594504F92402B5B5FADBDC0809120F9203928433DF1C14851DF461862AA2249";
    attribute INIT_29 of inst : label is "40100001100110011111100103351808000101B04094812AA8DD51C2082A3A79";
    attribute INIT_2A of inst : label is "0945028A040A2880048201020108250832020900004000000000050800144201";
    attribute INIT_2B of inst : label is "3A9197D51226DA8B08113AB344E2CD138B350C36D63003D83F926DB092000B05";
    attribute INIT_2C of inst : label is "4A9552859028FFD96651FFFFFF561896925922252900012AA2AA0A828051E93C";
    attribute INIT_2D of inst : label is "924924924924924924AAA853C12D2D1A4D14904BAD1A4D695429152AA952A800";
    attribute INIT_2E of inst : label is "0444812AA429142A74BA85481B656565CE72B2E7395957249249924924924924";
    attribute INIT_2F of inst : label is "FFFFFFFFFA88200A0A0A0A00A0003328D4600A0A288100847BA3B4B54D2DA0D1";
    attribute INIT_30 of inst : label is "1594504F92402B5B5FADBDC0809120F9203928433DF1C14851DF461862AA2249";
    attribute INIT_31 of inst : label is "40100001100110011111100103351808000101B04094812AA8DD51C2082A3A79";
    attribute INIT_32 of inst : label is "0945028A040A2880048201020108250832020900004000000000050800144201";
    attribute INIT_33 of inst : label is "3A9197D51226DA8B08113AB344E2CD138B350C36D63003D83F926DB092000B05";
    attribute INIT_34 of inst : label is "4A9552859028FFD96651FFFFFF561896925922252900012AA2AA0A828051E93C";
    attribute INIT_35 of inst : label is "924924924924924924AAA853C12D2D1A4D14904BAD1A4D695429152AA952A800";
    attribute INIT_36 of inst : label is "0444812AA429142A74BA85481B656565CE72B2E7395957249249924924924924";
    attribute INIT_37 of inst : label is "FFFFFFFFFA88200A0A0A0A00A0003328D4600A0A288100847BA3B4B54D2DA0D1";
    attribute INIT_38 of inst : label is "1594504F92402B5B5FADBDC0809120F9203928433DF1C14851DF461862AA2249";
    attribute INIT_39 of inst : label is "40100001100110011111100103351808000101B04094812AA8DD51C2082A3A79";
    attribute INIT_3A of inst : label is "0945028A040A2880048201020108250832020900004000000000050800144201";
    attribute INIT_3B of inst : label is "3A9197D51226DA8B08113AB344E2CD138B350C36D63003D83F926DB092000B05";
    attribute INIT_3C of inst : label is "4A9552859028FFD96651FFFFFF561896925922252900012AA2AA0A828051E93C";
    attribute INIT_3D of inst : label is "924924924924924924AAA853C12D2D1A4D14904BAD1A4D695429152AA952A800";
    attribute INIT_3E of inst : label is "0444812AA429142A74BA85481B656565CE72B2E7395957249249924924924924";
    attribute INIT_3F of inst : label is "FFFFFFFFFA88200A0A0A0A00A0003328D4600A0A288100847BA3B4B54D2DA0D1";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "06A2800008A2124D5F599BFCDCABBAC6F1076C21084BFF000000000000000000";
    attribute INIT_01 of inst : label is "FFFFFE3BFA009B7BFF1F048AC949AB591123FC1049A29A283C8B4C9706A10412";
    attribute INIT_02 of inst : label is "1A72C5864500D48A282D069B3B9A6C9334D926A9C02DB4F02B46AC61266C9ADF";
    attribute INIT_03 of inst : label is "5FFD898AFED206D2B423569B160387980D0F3122E36E356632BA1448746CFF60";
    attribute INIT_04 of inst : label is "F6812069269AB56AADAB56AAC2A0E197648B52926E9B29AD29D219C1AB709946";
    attribute INIT_05 of inst : label is "D12889415996C9249C90A92100C7116A305805B2E0891224482A4091109BFE5F";
    attribute INIT_06 of inst : label is "4A0AF44A04A04A44A4936E259C1F8A49B097B097B017B017B0DB914AD02C0780";
    attribute INIT_07 of inst : label is "1D830A0EC3AB0C8B0404A2EE63088A2D155892081208959040AC0828282B024A";
    attribute INIT_08 of inst : label is "494832E932EC836A529AD4A5FCDADA592D96CB6095095095095311A748560494";
    attribute INIT_09 of inst : label is "C8164A8B0888882A01104AC10474C460A17006C142F221845680D261B0890251";
    attribute INIT_0A of inst : label is "2949048160AD9648FFC11000BBE723C8430DC245F7908039130755555555F836";
    attribute INIT_0B of inst : label is "C033DD84400E96E02C09B6C9B6C9B6C9B6D42464B3C97C0276654B91BA187784";
    attribute INIT_0C of inst : label is "3009B4957218A89BCCBCE201B3C91240E62CC6A60C20136395112059895112C9";
    attribute INIT_0D of inst : label is "6FFFFFFFFF3573F85B593AD3B640A118888716FA87FC1C566D26B3C9FF1082DB";
    attribute INIT_0E of inst : label is "5480056A95AB00E820A96061960D39A1020C100D3A98C123D0294765B3650A37";
    attribute INIT_0F of inst : label is "0001FE7FF8003FC004000B00E71E236C4C4923B026C936409B24D9452900D985";
    attribute INIT_10 of inst : label is "06A2800008A2124D5F599BFCDCABBAC6F1076C21084BFF000000000000000000";
    attribute INIT_11 of inst : label is "FFFFFE3BFA009B7BFF1F048AC949AB591123FC1049A29A283C8B4C9706A10412";
    attribute INIT_12 of inst : label is "1A72C5864500D48A282D069B3B9A6C9334D926A9C02DB4F02B46AC61266C9ADF";
    attribute INIT_13 of inst : label is "5FFD898AFED206D2B423569B160387980D0F3122E36E356632BA1448746CFF60";
    attribute INIT_14 of inst : label is "F6812069269AB56AADAB56AAC2A0E197648B52926E9B29AD29D219C1AB709946";
    attribute INIT_15 of inst : label is "D12889415996C9249C90A92100C7116A305805B2E0891224482A4091109BFE5F";
    attribute INIT_16 of inst : label is "4A0AF44A04A04A44A4936E259C1F8A49B097B097B017B017B0DB914AD02C0780";
    attribute INIT_17 of inst : label is "1D830A0EC3AB0C8B0404A2EE63088A2D155892081208959040AC0828282B024A";
    attribute INIT_18 of inst : label is "494832E932EC836A529AD4A5FCDADA592D96CB6095095095095311A748560494";
    attribute INIT_19 of inst : label is "C8164A8B0888882A01104AC10474C460A17006C142F221845680D261B0890251";
    attribute INIT_1A of inst : label is "2949048160AD9648FFC11000BBE723C8430DC245F7908039130755555555F836";
    attribute INIT_1B of inst : label is "C033DD84400E96E02C09B6C9B6C9B6C9B6D42464B3C97C0276654B91BA187784";
    attribute INIT_1C of inst : label is "3009B4957218A89BCCBCE201B3C91240E62CC6A60C20136395112059895112C9";
    attribute INIT_1D of inst : label is "6FFFFFFFFF3573F85B593AD3B640A118888716FA87FC1C566D26B3C9FF1082DB";
    attribute INIT_1E of inst : label is "5480056A95AB00E820A96061960D39A1020C100D3A98C123D0294765B3650A37";
    attribute INIT_1F of inst : label is "0001FE7FF8003FC004000B00E71E236C4C4923B026C936409B24D9452900D985";
    attribute INIT_20 of inst : label is "31B3164C9249DA91C8F1783F83F200DB74DB2AD799BAC18C599B52B6F48AEA49";
    attribute INIT_21 of inst : label is "503303322223333220929AB90197030001010192421284271A4D5ADB613ADABB";
    attribute INIT_22 of inst : label is "0208041004104100450400040209275E26492492514400000000401C00065329";
    attribute INIT_23 of inst : label is "59C0482D7442D6B7998B6B826DAE09B698242026828002003F896CB249270088";
    attribute INIT_24 of inst : label is "BCE67D8B8B58FF42C0B7FFFFFF3E118DD1B5222B5916D958AB674A664CD6DD7B";
    attribute INIT_25 of inst : label is "924924924DA4D24924AA6A38E11514F399AC8C456AF399FCD3CE66D9A79CCC00";
    attribute INIT_26 of inst : label is "4E82DB59ABCE6669E7336CDDBD6565658C62B2C6315957349B49D24924924924";
    attribute INIT_27 of inst : label is "FFFFFFFFFFF7DFD76F7FFD5D5F4AF7B9946493830821103473336FA64BE921B8";
    attribute INIT_28 of inst : label is "31B3164C9249DA91C8F1783F83F200DB74DB2AD799BAC18C599B52B6F48AEA49";
    attribute INIT_29 of inst : label is "503303322223333220929AB90197030001010192421284271A4D5ADB613ADABB";
    attribute INIT_2A of inst : label is "0208041004104100450400040209275E26492492514400000000401C00065329";
    attribute INIT_2B of inst : label is "59C0482D7442D6B7998B6B826DAE09B698242026828002003F896CB249270088";
    attribute INIT_2C of inst : label is "BCE67D8B8B58FF42C0B7FFFFFF3E118DD1B5222B5916D958AB674A664CD6DD7B";
    attribute INIT_2D of inst : label is "924924924DA4D24924AA6A38E11514F399AC8C456AF399FCD3CE66D9A79CCC00";
    attribute INIT_2E of inst : label is "4E82DB59ABCE6669E7336CDDBD6565658C62B2C6315957349B49D24924924924";
    attribute INIT_2F of inst : label is "FFFFFFFFFFF7DFD76F7FFD5D5F4AF7B9946493830821103473336FA64BE921B8";
    attribute INIT_30 of inst : label is "31B3164C9249DA91C8F1783F83F200DB74DB2AD799BAC18C599B52B6F48AEA49";
    attribute INIT_31 of inst : label is "503303322223333220929AB90197030001010192421284271A4D5ADB613ADABB";
    attribute INIT_32 of inst : label is "0208041004104100450400040209275E26492492514400000000401C00065329";
    attribute INIT_33 of inst : label is "59C0482D7442D6B7998B6B826DAE09B698242026828002003F896CB249270088";
    attribute INIT_34 of inst : label is "BCE67D8B8B58FF42C0B7FFFFFF3E118DD1B5222B5916D958AB674A664CD6DD7B";
    attribute INIT_35 of inst : label is "924924924DA4D24924AA6A38E11514F399AC8C456AF399FCD3CE66D9A79CCC00";
    attribute INIT_36 of inst : label is "4E82DB59ABCE6669E7336CDDBD6565658C62B2C6315957349B49D24924924924";
    attribute INIT_37 of inst : label is "FFFFFFFFFFF7DFD76F7FFD5D5F4AF7B9946493830821103473336FA64BE921B8";
    attribute INIT_38 of inst : label is "31B3164C9249DA91C8F1783F83F200DB74DB2AD799BAC18C599B52B6F48AEA49";
    attribute INIT_39 of inst : label is "503303322223333220929AB90197030001010192421284271A4D5ADB613ADABB";
    attribute INIT_3A of inst : label is "0208041004104100450400040209275E26492492514400000000401C00065329";
    attribute INIT_3B of inst : label is "59C0482D7442D6B7998B6B826DAE09B698242026828002003F896CB249270088";
    attribute INIT_3C of inst : label is "BCE67D8B8B58FF42C0B7FFFFFF3E118DD1B5222B5916D958AB674A664CD6DD7B";
    attribute INIT_3D of inst : label is "924924924DA4D24924AA6A38E11514F399AC8C456AF399FCD3CE66D9A79CCC00";
    attribute INIT_3E of inst : label is "4E82DB59ABCE6669E7336CDDBD6565658C62B2C6315957349B49D24924924924";
    attribute INIT_3F of inst : label is "FFFFFFFFFFF7DFD76F7FFD5D5F4AF7B9946493830821103473336FA64BE921B8";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "F93CACCCF7F80938B764368C0C09EBDE6711F460917700000000000000000000";
    attribute INIT_01 of inst : label is "FFFFFF8622081AAE30313261242716B71107FED12E3CF3809E7632CC864C16DB";
    attribute INIT_02 of inst : label is "24C95331302E066184CB9450CB9A6C9334D926AE29D0912B969C5B8C3B1AF037";
    attribute INIT_03 of inst : label is "77FEEC3FA2461D80FB8C18E05C1E3C20787846859C11C1D9E8ED9B2F07D87F93";
    attribute INIT_04 of inst : label is "384C93049265CB97725CB9772381E443E0202459EA5EA1ACCFF03E261408F473";
    attribute INIT_05 of inst : label is "2CD96C6C7764A4920E5D14E2CB8103D3692C30419E74E9D3A4276ACDF0212419";
    attribute INIT_06 of inst : label is "2363035275275235234EC213044FE1656663A663A2E3A6E3A2A41623E49279CF";
    attribute INIT_07 of inst : label is "669D63334C8C770C04121E660CAF14DA44740165C92E4749723AED8D8D8CBB23";
    attribute INIT_08 of inst : label is "6D69C110C1000C841DE1083BFEB036361A0D068701F01F01F018D039831D76C6";
    attribute INIT_09 of inst : label is "3580306EDDB5DBD505DB239C0BC70B04128C8008252CA58146770B706406B90E";
    attribute INIT_0A of inst : label is "E52CB64D923B1240FFEFAAAAEEB22489A492F91F59130491049255555555FD80";
    attribute INIT_0B of inst : label is "FB608C0524780D04D0CF410741074107412CB39A6DB603F9CDD44665F8C87FB3";
    attribute INIT_0C of inst : label is "1B0D42C2C8726A6EE862385C4E25ED00F426335A163128D8ED4C232C64D4C274";
    attribute INIT_0D of inst : label is "0BFFFFFFFFC067FDAEA4E58E0D6E05C76E3D41BE04FEF52D90924822FFC6F1A4";
    attribute INIT_0E of inst : label is "B7001B96EE5C978DB22DD31F4392650D6D965992616CE68FEC849CDC7A4201A8";
    attribute INIT_0F of inst : label is "0001027FF800204004032610B2E43C813AC61C4BB605B02ED816C07185C9EC70";
    attribute INIT_10 of inst : label is "F93CACCCF7F80938B764368C0C09EBDE6711F460917700000000000000000000";
    attribute INIT_11 of inst : label is "FFFFFF8622081AAE30313261242716B71107FED12E3CF3809E7632CC864C16DB";
    attribute INIT_12 of inst : label is "24C95331302E066184CB9450CB9A6C9334D926AE29D0912B969C5B8C3B1AF037";
    attribute INIT_13 of inst : label is "77FEEC3FA2461D80FB8C18E05C1E3C20787846859C11C1D9E8ED9B2F07D87F93";
    attribute INIT_14 of inst : label is "384C93049265CB97725CB9772381E443E0202459EA5EA1ACCFF03E261408F473";
    attribute INIT_15 of inst : label is "2CD96C6C7764A4920E5D14E2CB8103D3692C30419E74E9D3A4276ACDF0212419";
    attribute INIT_16 of inst : label is "2363035275275235234EC213044FE1656663A663A2E3A6E3A2A41623E49279CF";
    attribute INIT_17 of inst : label is "669D63334C8C770C04121E660CAF14DA44740165C92E4749723AED8D8D8CBB23";
    attribute INIT_18 of inst : label is "6D69C110C1000C841DE1083BFEB036361A0D068701F01F01F018D039831D76C6";
    attribute INIT_19 of inst : label is "3580306EDDB5DBD505DB239C0BC70B04128C8008252CA58146770B706406B90E";
    attribute INIT_1A of inst : label is "E52CB64D923B1240FFEFAAAAEEB22489A492F91F59130491049255555555FD80";
    attribute INIT_1B of inst : label is "FB608C0524780D04D0CF410741074107412CB39A6DB603F9CDD44665F8C87FB3";
    attribute INIT_1C of inst : label is "1B0D42C2C8726A6EE862385C4E25ED00F426335A163128D8ED4C232C64D4C274";
    attribute INIT_1D of inst : label is "0BFFFFFFFFC067FDAEA4E58E0D6E05C76E3D41BE04FEF52D90924822FFC6F1A4";
    attribute INIT_1E of inst : label is "B7001B96EE5C978DB22DD31F4392650D6D965992616CE68FEC849CDC7A4201A8";
    attribute INIT_1F of inst : label is "0001027FF800204004032610B2E43C813AC61C4BB605B02ED816C07185C9EC70";
    attribute INIT_20 of inst : label is "9CD9E13ACB30FB5B5AFD38A28459B396C2158DA84324A56B643229418760232C";
    attribute INIT_21 of inst : label is "501111111110000001C1C00C009505010101019598493092D52824B4CDCD912D";
    attribute INIT_22 of inst : label is "6C92592497649249724925CB259490B19909249240400000000045044147000C";
    attribute INIT_23 of inst : label is "951FF6C88BBD840526E36A938DAA4E36A93244B8C81093487FC9FB0849249092";
    attribute INIT_24 of inst : label is "61088132E691FF249921FFFFFFA32C692C21989294C006960054A341386C921A";
    attribute INIT_25 of inst : label is "9249A4924924924926AB438C01C9C384224AE2704184227E8E1088151C211240";
    attribute INIT_26 of inst : label is "B9370495061089C708441AB04B6565656B5AB2B5AD595726D2491A4924924D24";
    attribute INIT_27 of inst : label is "FFFFFFFFF88AAA888022200A2E242A2CE35268C866DE48C7BC82E49109348491";
    attribute INIT_28 of inst : label is "9CD9E13ACB30FB5B5AFD38A28459B396C2158DA84324A56B643229418760232C";
    attribute INIT_29 of inst : label is "501111111110000001C1C00C009505010101019598493092D52824B4CDCD912D";
    attribute INIT_2A of inst : label is "6C92592497649249724925CB259490B19909249240400000000045044147000C";
    attribute INIT_2B of inst : label is "951FF6C88BBD840526E36A938DAA4E36A93244B8C81093487FC9FB0849249092";
    attribute INIT_2C of inst : label is "61088132E691FF249921FFFFFFA32C692C21989294C006960054A341386C921A";
    attribute INIT_2D of inst : label is "9249A4924924924926AB438C01C9C384224AE2704184227E8E1088151C211240";
    attribute INIT_2E of inst : label is "B9370495061089C708441AB04B6565656B5AB2B5AD595726D2491A4924924D24";
    attribute INIT_2F of inst : label is "FFFFFFFFF88AAA888022200A2E242A2CE35268C866DE48C7BC82E49109348491";
    attribute INIT_30 of inst : label is "9CD9E13ACB30FB5B5AFD38A28459B396C2158DA84324A56B643229418760232C";
    attribute INIT_31 of inst : label is "501111111110000001C1C00C009505010101019598493092D52824B4CDCD912D";
    attribute INIT_32 of inst : label is "6C92592497649249724925CB259490B19909249240400000000045044147000C";
    attribute INIT_33 of inst : label is "951FF6C88BBD840526E36A938DAA4E36A93244B8C81093487FC9FB0849249092";
    attribute INIT_34 of inst : label is "61088132E691FF249921FFFFFFA32C692C21989294C006960054A341386C921A";
    attribute INIT_35 of inst : label is "9249A4924924924926AB438C01C9C384224AE2704184227E8E1088151C211240";
    attribute INIT_36 of inst : label is "B9370495061089C708441AB04B6565656B5AB2B5AD595726D2491A4924924D24";
    attribute INIT_37 of inst : label is "FFFFFFFFF88AAA888022200A2E242A2CE35268C866DE48C7BC82E49109348491";
    attribute INIT_38 of inst : label is "9CD9E13ACB30FB5B5AFD38A28459B396C2158DA84324A56B643229418760232C";
    attribute INIT_39 of inst : label is "501111111110000001C1C00C009505010101019598493092D52824B4CDCD912D";
    attribute INIT_3A of inst : label is "6C92592497649249724925CB259490B19909249240400000000045044147000C";
    attribute INIT_3B of inst : label is "951FF6C88BBD840526E36A938DAA4E36A93244B8C81093487FC9FB0849249092";
    attribute INIT_3C of inst : label is "61088132E691FF249921FFFFFFA32C692C21989294C006960054A341386C921A";
    attribute INIT_3D of inst : label is "9249A4924924924926AB438C01C9C384224AE2704184227E8E1088151C211240";
    attribute INIT_3E of inst : label is "B9370495061089C708441AB04B6565656B5AB2B5AD595726D2491A4924924D24";
    attribute INIT_3F of inst : label is "FFFFFFFFF88AAA888022200A2E242A2CE35268C866DE48C7BC82E49109348491";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "F155BDDDD7F80DA8D7AC62040C19A74E670BFC24205700000000000000000000";
    attribute INIT_01 of inst : label is "FFFFFF86A002BE0C21320940A2B51AD60007FF533451455197D2128487D81FED";
    attribute INIT_02 of inst : label is "1450217228B5445146FBFC71AD534ADAA695B4AD6B0000091AB46A88592AD057";
    attribute INIT_03 of inst : label is "57FEE83C80061481FFC88050542AD600A8AC0B1E8A28A151A8AC9B6603487FDB";
    attribute INIT_04 of inst : label is "2158D630C3408102200810222301A223E196A151E35B856E8EE03D651A18D4E3";
    attribute INIT_05 of inst : label is "A4893474552D80000F6F18EA6B42036B2BEC6220A3468D1A3437B24DF0000010";
    attribute INIT_06 of inst : label is "E3E20F18B18B18B18B80C003000FD14726E3626362E3666363929627E78BF5FE";
    attribute INIT_07 of inst : label is "C775E3E3B888514000121E6708A404EA445641B48FFEC57FF62BEF8F8F88FBE3";
    attribute INIT_08 of inst : label is "6F7FA8BCA8A60A4728D08E51FF90541A0C06030542D42D42D42AD4D1E715F7C7";
    attribute INIT_09 of inst : label is "17C311EA88F08F8007DDA288095289367347926CE6ADB503CC7E8B51660ADD3B";
    attribute INIT_0A of inst : label is "E73EFB6D9A2B0018FFD44555C00A0280A288F46805010450028A00000000FFC3";
    attribute INIT_0B of inst : label is "C9608C8C346A14BFE9D5829D829D829D82849F59018680035554426DF0887F93";
    attribute INIT_0C of inst : label is "1D1F228A41702032F80635EADC66A600F4063A0C1C71A050C4080A2C70408060";
    attribute INIT_0D of inst : label is "3BFFFFFFFFA05FFEB2D7AEBA95FD1E87F47482BE06FFD23500020006FF8BF292";
    attribute INIT_0E of inst : label is "280011034408FEA79E255A1D238A2F1D3C934F8A2F6CF717E4421CDCBEC327E8";
    attribute INIT_0F of inst : label is "000100000800004000013604B2D05A41EC62780FB465A33ED1968C210EEFEC62";
    attribute INIT_10 of inst : label is "F155BDDDD7F80DA8D7AC62040C19A74E670BFC24205700000000000000000000";
    attribute INIT_11 of inst : label is "FFFFFF86A002BE0C21320940A2B51AD60007FF533451455197D2128487D81FED";
    attribute INIT_12 of inst : label is "1450217228B5445146FBFC71AD534ADAA695B4AD6B0000091AB46A88592AD057";
    attribute INIT_13 of inst : label is "57FEE83C80061481FFC88050542AD600A8AC0B1E8A28A151A8AC9B6603487FDB";
    attribute INIT_14 of inst : label is "2158D630C3408102200810222301A223E196A151E35B856E8EE03D651A18D4E3";
    attribute INIT_15 of inst : label is "A4893474552D80000F6F18EA6B42036B2BEC6220A3468D1A3437B24DF0000010";
    attribute INIT_16 of inst : label is "E3E20F18B18B18B18B80C003000FD14726E3626362E3666363929627E78BF5FE";
    attribute INIT_17 of inst : label is "C775E3E3B888514000121E6708A404EA445641B48FFEC57FF62BEF8F8F88FBE3";
    attribute INIT_18 of inst : label is "6F7FA8BCA8A60A4728D08E51FF90541A0C06030542D42D42D42AD4D1E715F7C7";
    attribute INIT_19 of inst : label is "17C311EA88F08F8007DDA288095289367347926CE6ADB503CC7E8B51660ADD3B";
    attribute INIT_1A of inst : label is "E73EFB6D9A2B0018FFD44555C00A0280A288F46805010450028A00000000FFC3";
    attribute INIT_1B of inst : label is "C9608C8C346A14BFE9D5829D829D829D82849F59018680035554426DF0887F93";
    attribute INIT_1C of inst : label is "1D1F228A41702032F80635EADC66A600F4063A0C1C71A050C4080A2C70408060";
    attribute INIT_1D of inst : label is "3BFFFFFFFFA05FFEB2D7AEBA95FD1E87F47482BE06FFD23500020006FF8BF292";
    attribute INIT_1E of inst : label is "280011034408FEA79E255A1D238A2F1D3C934F8A2F6CF717E4421CDCBEC327E8";
    attribute INIT_1F of inst : label is "000100000800004000013604B2D05A41EC62780FB465A33ED1968C210EEFEC62";
    attribute INIT_20 of inst : label is "88F882028A30F9494AFA30630211DEB25E778EB4C66FBDED6C6631A285502228";
    attribute INIT_21 of inst : label is "103323333333333332828AF8009C06040000008CB1C5638BF63897905480B1EF";
    attribute INIT_22 of inst : label is "779E6F3CBFBCF3CBFBCF2FD92C9003C388092492510000000000451401521428";
    attribute INIT_23 of inst : label is "F76C46D8EDB48C1DFED1288944A2251288920314480F6947BFC9E1004925B0BE";
    attribute INIT_24 of inst : label is "3008077EC0F7FF6799E2FFFFFFEB643B64E1111EF08042F501DDC1C02805B616";
    attribute INIT_25 of inst : label is "DB6DB6DB6DB6DB6DB6ABC51800A8A2C0207B5428C0C020778B008077160103C0";
    attribute INIT_26 of inst : label is "AB220AF70300814580402B94AD15151508428A84214556B6DB6D5B6DB6DB6DB6";
    attribute INIT_27 of inst : label is "FFFFFFFFFA220EA8A28282202F9422F2A24920C0441F085A9412640209000088";
    attribute INIT_28 of inst : label is "88F882028A30F9494AFA30630211DEB25E778EB4C66FBDED6C6631A285502228";
    attribute INIT_29 of inst : label is "103323333333333332828AF8009C06040000008CB1C5638BF63897905480B1EF";
    attribute INIT_2A of inst : label is "779E6F3CBFBCF3CBFBCF2FD92C9003C388092492510000000000451401521428";
    attribute INIT_2B of inst : label is "F76C46D8EDB48C1DFED1288944A2251288920314480F6947BFC9E1004925B0BE";
    attribute INIT_2C of inst : label is "3008077EC0F7FF6799E2FFFFFFEB643B64E1111EF08042F501DDC1C02805B616";
    attribute INIT_2D of inst : label is "DB6DB6DB6DB6DB6DB6ABC51800A8A2C0207B5428C0C020778B008077160103C0";
    attribute INIT_2E of inst : label is "AB220AF70300814580402B94AD15151508428A84214556B6DB6D5B6DB6DB6DB6";
    attribute INIT_2F of inst : label is "FFFFFFFFFA220EA8A28282202F9422F2A24920C0441F085A9412640209000088";
    attribute INIT_30 of inst : label is "88F882028A30F9494AFA30630211DEB25E778EB4C66FBDED6C6631A285502228";
    attribute INIT_31 of inst : label is "103323333333333332828AF8009C06040000008CB1C5638BF63897905480B1EF";
    attribute INIT_32 of inst : label is "779E6F3CBFBCF3CBFBCF2FD92C9003C388092492510000000000451401521428";
    attribute INIT_33 of inst : label is "F76C46D8EDB48C1DFED1288944A2251288920314480F6947BFC9E1004925B0BE";
    attribute INIT_34 of inst : label is "3008077EC0F7FF6799E2FFFFFFEB643B64E1111EF08042F501DDC1C02805B616";
    attribute INIT_35 of inst : label is "DB6DB6DB6DB6DB6DB6ABC51800A8A2C0207B5428C0C020778B008077160103C0";
    attribute INIT_36 of inst : label is "AB220AF70300814580402B94AD15151508428A84214556B6DB6D5B6DB6DB6DB6";
    attribute INIT_37 of inst : label is "FFFFFFFFFA220EA8A28282202F9422F2A24920C0441F085A9412640209000088";
    attribute INIT_38 of inst : label is "88F882028A30F9494AFA30630211DEB25E778EB4C66FBDED6C6631A285502228";
    attribute INIT_39 of inst : label is "103323333333333332828AF8009C06040000008CB1C5638BF63897905480B1EF";
    attribute INIT_3A of inst : label is "779E6F3CBFBCF3CBFBCF2FD92C9003C388092492510000000000451401521428";
    attribute INIT_3B of inst : label is "F76C46D8EDB48C1DFED1288944A2251288920314480F6947BFC9E1004925B0BE";
    attribute INIT_3C of inst : label is "3008077EC0F7FF6799E2FFFFFFEB643B64E1111EF08042F501DDC1C02805B616";
    attribute INIT_3D of inst : label is "DB6DB6DB6DB6DB6DB6ABC51800A8A2C0207B5428C0C020778B008077160103C0";
    attribute INIT_3E of inst : label is "AB220AF70300814580402B94AD15151508428A84214556B6DB6D5B6DB6DB6DB6";
    attribute INIT_3F of inst : label is "FFFFFFFFFA220EA8A28282202F9422F2A24920C0441F085A9412640209000088";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
