library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sprom_jiffy is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sprom_jiffy is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"97",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"78",X"A9",X"F7",X"2D",X"00",X"1C",X"48",X"A5",X"7F",X"F0",X"05",X"68",X"09",X"00",X"D0",X"03",
		X"68",X"09",X"08",X"8D",X"00",X"1C",X"58",X"60",X"78",X"A9",X"08",X"0D",X"00",X"1C",X"8D",X"00",
		X"1C",X"58",X"60",X"A9",X"00",X"8D",X"6C",X"02",X"8D",X"6D",X"02",X"60",X"78",X"8A",X"48",X"A9",
		X"50",X"8D",X"6C",X"02",X"A2",X"00",X"BD",X"CA",X"FE",X"8D",X"6D",X"02",X"0D",X"00",X"1C",X"8D",
		X"00",X"1C",X"68",X"AA",X"58",X"60",X"A9",X"00",X"8D",X"F9",X"02",X"AD",X"8E",X"02",X"85",X"7F",
		X"20",X"BC",X"E6",X"A5",X"84",X"10",X"09",X"29",X"0F",X"C9",X"0F",X"F0",X"03",X"4C",X"B4",X"D7",
		X"20",X"B3",X"C2",X"B1",X"A3",X"8D",X"75",X"02",X"A2",X"0B",X"BD",X"89",X"FE",X"CD",X"75",X"02",
		X"F0",X"08",X"CA",X"10",X"F5",X"A9",X"31",X"4C",X"C8",X"C1",X"8E",X"2A",X"02",X"E0",X"09",X"90",
		X"03",X"20",X"EE",X"C1",X"AE",X"2A",X"02",X"BD",X"95",X"FE",X"85",X"6F",X"BD",X"A1",X"FE",X"85",
		X"70",X"6C",X"6F",X"00",X"A9",X"00",X"8D",X"F9",X"02",X"AD",X"6C",X"02",X"D0",X"2A",X"A0",X"00",
		X"98",X"84",X"80",X"84",X"81",X"84",X"A3",X"20",X"C7",X"E6",X"20",X"23",X"C1",X"A5",X"7F",X"8D",
		X"8E",X"02",X"AA",X"A9",X"00",X"95",X"FF",X"20",X"BD",X"C1",X"4C",X"DA",X"D4",X"A0",X"28",X"A9",
		X"00",X"99",X"00",X"02",X"88",X"10",X"FA",X"60",X"A0",X"00",X"84",X"80",X"84",X"81",X"4C",X"45",
		X"E6",X"A2",X"00",X"8E",X"7A",X"02",X"A9",X"3A",X"20",X"68",X"C2",X"F0",X"05",X"88",X"88",X"8C",
		X"7A",X"02",X"4C",X"68",X"C3",X"A0",X"00",X"A2",X"00",X"A9",X"3A",X"4C",X"68",X"C2",X"20",X"E5",
		X"C1",X"D0",X"05",X"A9",X"34",X"4C",X"C8",X"C1",X"88",X"88",X"8C",X"7A",X"02",X"8A",X"D0",X"F3",
		X"A9",X"3D",X"20",X"68",X"C2",X"8A",X"F0",X"02",X"A9",X"40",X"09",X"21",X"8D",X"8B",X"02",X"E8",
		X"8E",X"77",X"02",X"8E",X"78",X"02",X"AD",X"8A",X"02",X"F0",X"0D",X"A9",X"80",X"0D",X"8B",X"02",
		X"8D",X"8B",X"02",X"A9",X"00",X"8D",X"8A",X"02",X"98",X"F0",X"29",X"9D",X"7A",X"02",X"AD",X"77",
		X"02",X"8D",X"79",X"02",X"A9",X"8D",X"20",X"68",X"C2",X"E8",X"8E",X"78",X"02",X"CA",X"AD",X"8A",
		X"02",X"F0",X"02",X"A9",X"08",X"EC",X"77",X"02",X"F0",X"02",X"09",X"04",X"09",X"03",X"4D",X"8B",
		X"02",X"8D",X"8B",X"02",X"AD",X"8B",X"02",X"AE",X"2A",X"02",X"3D",X"A5",X"FE",X"D0",X"01",X"60",
		X"8D",X"6C",X"02",X"A9",X"30",X"4C",X"C8",X"C1",X"8D",X"75",X"02",X"CC",X"74",X"02",X"B0",X"2E",
		X"B1",X"A3",X"C8",X"CD",X"75",X"02",X"F0",X"28",X"C9",X"2A",X"F0",X"04",X"C9",X"3F",X"D0",X"03",
		X"EE",X"8A",X"02",X"C9",X"2C",X"D0",X"E4",X"98",X"9D",X"7B",X"02",X"AD",X"8A",X"02",X"29",X"7F",
		X"F0",X"07",X"A9",X"80",X"95",X"E7",X"8D",X"8A",X"02",X"E8",X"E0",X"04",X"90",X"CD",X"A0",X"00",
		X"AD",X"74",X"02",X"9D",X"7B",X"02",X"AD",X"8A",X"02",X"29",X"7F",X"F0",X"04",X"A9",X"80",X"95",
		X"E7",X"98",X"60",X"A4",X"A3",X"F0",X"14",X"88",X"F0",X"10",X"B9",X"00",X"02",X"C9",X"0D",X"F0",
		X"0A",X"88",X"B9",X"00",X"02",X"C9",X"0D",X"F0",X"02",X"C8",X"C8",X"8C",X"74",X"02",X"C0",X"2A",
		X"A0",X"FF",X"90",X"08",X"8C",X"2A",X"02",X"A9",X"32",X"4C",X"C8",X"C1",X"A0",X"00",X"98",X"85",
		X"A3",X"8D",X"58",X"02",X"8D",X"4A",X"02",X"8D",X"96",X"02",X"85",X"D3",X"8D",X"79",X"02",X"8D",
		X"77",X"02",X"8D",X"78",X"02",X"8D",X"8A",X"02",X"8D",X"6C",X"02",X"A2",X"05",X"9D",X"79",X"02",
		X"95",X"D7",X"95",X"DC",X"95",X"E1",X"95",X"E6",X"9D",X"7F",X"02",X"9D",X"84",X"02",X"CA",X"D0",
		X"EC",X"60",X"AD",X"78",X"02",X"8D",X"77",X"02",X"A9",X"01",X"8D",X"78",X"02",X"8D",X"79",X"02",
		X"AC",X"8E",X"02",X"A2",X"00",X"86",X"D3",X"BD",X"7A",X"02",X"20",X"3C",X"C3",X"A6",X"D3",X"9D",
		X"7A",X"02",X"98",X"95",X"E2",X"E8",X"EC",X"78",X"02",X"90",X"EA",X"60",X"AA",X"A0",X"00",X"A9",
		X"3A",X"DD",X"01",X"02",X"F0",X"0C",X"DD",X"00",X"02",X"D0",X"16",X"E8",X"98",X"29",X"01",X"A8",
		X"8A",X"60",X"BD",X"00",X"02",X"E8",X"E8",X"C9",X"30",X"F0",X"F2",X"C9",X"31",X"F0",X"EE",X"D0",
		X"EB",X"98",X"09",X"80",X"29",X"81",X"D0",X"E7",X"A9",X"00",X"8D",X"8B",X"02",X"AC",X"7A",X"02",
		X"B1",X"A3",X"20",X"BD",X"C3",X"10",X"11",X"C8",X"CC",X"74",X"02",X"B0",X"06",X"AC",X"74",X"02",
		X"88",X"D0",X"ED",X"CE",X"8B",X"02",X"A9",X"00",X"29",X"01",X"85",X"7F",X"4C",X"00",X"C1",X"A5",
		X"7F",X"49",X"01",X"29",X"01",X"85",X"7F",X"60",X"A0",X"00",X"AD",X"77",X"02",X"CD",X"78",X"02",
		X"F0",X"16",X"CE",X"78",X"02",X"AC",X"78",X"02",X"B9",X"7A",X"02",X"A8",X"B1",X"A3",X"A0",X"04",
		X"D9",X"BB",X"FE",X"F0",X"03",X"88",X"D0",X"F8",X"98",X"8D",X"96",X"02",X"60",X"C9",X"30",X"F0",
		X"06",X"C9",X"31",X"F0",X"02",X"09",X"80",X"29",X"81",X"60",X"A9",X"00",X"85",X"6F",X"8D",X"8D",
		X"02",X"48",X"AE",X"78",X"02",X"68",X"05",X"6F",X"48",X"A9",X"01",X"85",X"6F",X"CA",X"30",X"0F",
		X"B5",X"E2",X"10",X"04",X"06",X"6F",X"06",X"6F",X"4A",X"90",X"EA",X"06",X"6F",X"D0",X"E6",X"68",
		X"AA",X"BD",X"3F",X"C4",X"48",X"29",X"03",X"8D",X"8C",X"02",X"68",X"0A",X"10",X"3E",X"A5",X"E2",
		X"29",X"01",X"85",X"7F",X"AD",X"8C",X"02",X"F0",X"2B",X"20",X"3D",X"C6",X"F0",X"12",X"20",X"8F",
		X"C3",X"A9",X"00",X"8D",X"8C",X"02",X"20",X"3D",X"C6",X"F0",X"1E",X"A9",X"74",X"20",X"C8",X"C1",
		X"20",X"8F",X"C3",X"20",X"3D",X"C6",X"08",X"20",X"8F",X"C3",X"28",X"F0",X"0C",X"A9",X"00",X"8D",
		X"8C",X"02",X"F0",X"05",X"20",X"3D",X"C6",X"D0",X"E2",X"4C",X"00",X"C1",X"2A",X"4C",X"00",X"C4",
		X"00",X"80",X"41",X"01",X"01",X"01",X"01",X"81",X"81",X"81",X"81",X"42",X"42",X"42",X"42",X"20",
		X"CA",X"C3",X"A9",X"00",X"8D",X"92",X"02",X"20",X"AC",X"C5",X"D0",X"19",X"CE",X"8C",X"02",X"10",
		X"01",X"60",X"A9",X"01",X"8D",X"8D",X"02",X"20",X"8F",X"C3",X"20",X"00",X"C1",X"4C",X"52",X"C4",
		X"20",X"17",X"C6",X"F0",X"10",X"20",X"D8",X"C4",X"AD",X"8F",X"02",X"F0",X"01",X"60",X"AD",X"53",
		X"02",X"30",X"ED",X"10",X"F0",X"AD",X"8F",X"02",X"F0",X"D2",X"60",X"20",X"04",X"C6",X"F0",X"1A",
		X"D0",X"28",X"A9",X"01",X"8D",X"8D",X"02",X"20",X"8F",X"C3",X"20",X"00",X"C1",X"A9",X"00",X"8D",
		X"92",X"02",X"20",X"AC",X"C5",X"D0",X"13",X"8D",X"8F",X"02",X"AD",X"8F",X"02",X"D0",X"28",X"CE",
		X"8C",X"02",X"10",X"DE",X"60",X"20",X"17",X"C6",X"F0",X"F0",X"20",X"D8",X"C4",X"AE",X"53",X"02",
		X"10",X"07",X"AD",X"8F",X"02",X"F0",X"EE",X"D0",X"0E",X"AD",X"96",X"02",X"F0",X"09",X"B5",X"E7",
		X"29",X"07",X"CD",X"96",X"02",X"D0",X"DE",X"60",X"A2",X"FF",X"8E",X"53",X"02",X"E8",X"8E",X"8A",
		X"02",X"20",X"89",X"C5",X"F0",X"06",X"60",X"20",X"94",X"C5",X"D0",X"FA",X"A5",X"7F",X"55",X"E2",
		X"4A",X"90",X"0B",X"29",X"40",X"F0",X"F0",X"A9",X"02",X"CD",X"8C",X"02",X"F0",X"E9",X"BD",X"7A",
		X"02",X"AA",X"20",X"A6",X"C6",X"A0",X"03",X"4C",X"1D",X"C5",X"BD",X"00",X"02",X"D1",X"94",X"F0",
		X"0A",X"C9",X"3F",X"D0",X"D2",X"B1",X"94",X"C9",X"A0",X"F0",X"CC",X"E8",X"C8",X"EC",X"76",X"02",
		X"B0",X"09",X"BD",X"00",X"02",X"C9",X"2A",X"F0",X"0C",X"D0",X"DF",X"C0",X"13",X"B0",X"06",X"B1",
		X"94",X"C9",X"A0",X"D0",X"B2",X"AE",X"79",X"02",X"8E",X"53",X"02",X"B5",X"E7",X"29",X"80",X"8D",
		X"8A",X"02",X"AD",X"94",X"02",X"95",X"DD",X"A5",X"81",X"95",X"D8",X"A0",X"00",X"B1",X"94",X"C8",
		X"48",X"29",X"40",X"85",X"6F",X"68",X"29",X"DF",X"30",X"02",X"09",X"20",X"29",X"27",X"05",X"6F",
		X"85",X"6F",X"A9",X"80",X"35",X"E7",X"05",X"6F",X"95",X"E7",X"B5",X"E2",X"29",X"80",X"05",X"7F",
		X"95",X"E2",X"B1",X"94",X"9D",X"80",X"02",X"C8",X"B1",X"94",X"9D",X"85",X"02",X"AD",X"58",X"02",
		X"D0",X"07",X"A0",X"15",X"B1",X"94",X"8D",X"58",X"02",X"A9",X"FF",X"8D",X"8F",X"02",X"AD",X"78",
		X"02",X"8D",X"79",X"02",X"CE",X"79",X"02",X"10",X"01",X"60",X"AE",X"79",X"02",X"B5",X"E7",X"30",
		X"05",X"BD",X"80",X"02",X"D0",X"EE",X"A9",X"00",X"8D",X"8F",X"02",X"60",X"A0",X"00",X"8C",X"91",
		X"02",X"88",X"8C",X"53",X"02",X"AD",X"85",X"FE",X"85",X"80",X"A9",X"01",X"85",X"81",X"8D",X"93",
		X"02",X"20",X"75",X"D4",X"AD",X"93",X"02",X"D0",X"01",X"60",X"A9",X"07",X"8D",X"95",X"02",X"A9",
		X"00",X"20",X"F6",X"D4",X"8D",X"93",X"02",X"20",X"E8",X"D4",X"CE",X"95",X"02",X"A0",X"00",X"B1",
		X"94",X"D0",X"18",X"AD",X"91",X"02",X"D0",X"2F",X"20",X"3B",X"DE",X"A5",X"81",X"8D",X"91",X"02",
		X"A5",X"94",X"AE",X"92",X"02",X"8D",X"92",X"02",X"F0",X"1D",X"60",X"A2",X"01",X"EC",X"92",X"02",
		X"D0",X"2D",X"F0",X"13",X"AD",X"85",X"FE",X"85",X"80",X"AD",X"90",X"02",X"85",X"81",X"20",X"75",
		X"D4",X"AD",X"94",X"02",X"20",X"C8",X"D4",X"A9",X"FF",X"8D",X"53",X"02",X"AD",X"95",X"02",X"30",
		X"08",X"A9",X"20",X"20",X"C6",X"D1",X"4C",X"D7",X"C5",X"20",X"4D",X"D4",X"4C",X"C4",X"C5",X"A5",
		X"94",X"8D",X"94",X"02",X"20",X"3B",X"DE",X"A5",X"81",X"8D",X"90",X"02",X"60",X"A5",X"68",X"D0",
		X"28",X"A6",X"7F",X"56",X"1C",X"90",X"22",X"A9",X"FF",X"8D",X"98",X"02",X"20",X"0E",X"D0",X"A0",
		X"FF",X"C9",X"02",X"F0",X"0A",X"C9",X"03",X"F0",X"06",X"C9",X"0F",X"F0",X"02",X"A0",X"00",X"A6",
		X"7F",X"98",X"95",X"FF",X"D0",X"03",X"20",X"42",X"D0",X"A6",X"7F",X"B5",X"FF",X"60",X"48",X"20",
		X"A6",X"C6",X"20",X"88",X"C6",X"68",X"38",X"ED",X"4B",X"02",X"AA",X"F0",X"0A",X"90",X"08",X"A9",
		X"A0",X"91",X"94",X"C8",X"CA",X"D0",X"FA",X"60",X"98",X"0A",X"A8",X"B9",X"99",X"00",X"85",X"94",
		X"B9",X"9A",X"00",X"85",X"95",X"A0",X"00",X"BD",X"00",X"02",X"91",X"94",X"C8",X"F0",X"06",X"E8",
		X"EC",X"76",X"02",X"90",X"F2",X"60",X"A9",X"00",X"8D",X"4B",X"02",X"8A",X"48",X"BD",X"00",X"02",
		X"C9",X"2C",X"F0",X"14",X"C9",X"3D",X"F0",X"10",X"EE",X"4B",X"02",X"E8",X"A9",X"0F",X"CD",X"4B",
		X"02",X"90",X"05",X"EC",X"74",X"02",X"90",X"E5",X"8E",X"76",X"02",X"68",X"AA",X"60",X"A5",X"83",
		X"48",X"A5",X"82",X"48",X"20",X"DE",X"C6",X"68",X"85",X"82",X"68",X"85",X"83",X"60",X"A9",X"11",
		X"85",X"83",X"20",X"EB",X"D0",X"20",X"E8",X"D4",X"AD",X"53",X"02",X"10",X"0A",X"AD",X"8D",X"02",
		X"D0",X"0A",X"20",X"06",X"C8",X"18",X"60",X"AD",X"8D",X"02",X"F0",X"1F",X"CE",X"8D",X"02",X"D0",
		X"0D",X"CE",X"8D",X"02",X"20",X"8F",X"C3",X"20",X"06",X"C8",X"38",X"4C",X"8F",X"C3",X"A9",X"00",
		X"8D",X"73",X"02",X"8D",X"8D",X"02",X"20",X"B7",X"C7",X"38",X"60",X"A2",X"18",X"A0",X"1D",X"B1",
		X"94",X"8D",X"73",X"02",X"F0",X"02",X"A2",X"16",X"88",X"B1",X"94",X"8D",X"72",X"02",X"E0",X"16",
		X"F0",X"0A",X"C9",X"0A",X"90",X"06",X"CA",X"C9",X"64",X"90",X"01",X"CA",X"20",X"AC",X"C7",X"B1",
		X"94",X"48",X"0A",X"10",X"05",X"A9",X"3C",X"9D",X"B2",X"02",X"68",X"29",X"0F",X"A8",X"B9",X"C5",
		X"FE",X"9D",X"B1",X"02",X"CA",X"B9",X"C0",X"FE",X"9D",X"B1",X"02",X"CA",X"B9",X"BB",X"FE",X"9D",
		X"B1",X"02",X"CA",X"CA",X"B0",X"05",X"A9",X"2A",X"9D",X"B2",X"02",X"A9",X"A0",X"9D",X"B1",X"02",
		X"CA",X"A0",X"12",X"B1",X"94",X"9D",X"B1",X"02",X"CA",X"88",X"C0",X"03",X"B0",X"F5",X"A9",X"22",
		X"9D",X"B1",X"02",X"E8",X"E0",X"20",X"B0",X"0B",X"BD",X"B1",X"02",X"C9",X"22",X"F0",X"04",X"C9",
		X"A0",X"D0",X"F0",X"A9",X"22",X"9D",X"B1",X"02",X"E8",X"E0",X"20",X"B0",X"0A",X"A9",X"7F",X"3D",
		X"B1",X"02",X"9D",X"B1",X"02",X"10",X"F1",X"20",X"B5",X"C4",X"38",X"60",X"A0",X"1B",X"A9",X"20",
		X"99",X"B0",X"02",X"88",X"D0",X"FA",X"60",X"20",X"19",X"F1",X"20",X"DF",X"F0",X"20",X"AC",X"C7",
		X"A9",X"FF",X"85",X"6F",X"A6",X"7F",X"8E",X"72",X"02",X"A9",X"00",X"8D",X"73",X"02",X"A6",X"F9",
		X"BD",X"E0",X"FE",X"85",X"95",X"AD",X"88",X"FE",X"85",X"94",X"A0",X"16",X"B1",X"94",X"C9",X"A0",
		X"D0",X"0B",X"A9",X"31",X"2C",X"B1",X"94",X"C9",X"A0",X"D0",X"02",X"A9",X"20",X"99",X"B3",X"02",
		X"88",X"10",X"F2",X"A9",X"12",X"8D",X"B1",X"02",X"A9",X"22",X"8D",X"B2",X"02",X"8D",X"C3",X"02",
		X"A9",X"20",X"8D",X"C4",X"02",X"60",X"20",X"AC",X"C7",X"A0",X"0B",X"B9",X"17",X"C8",X"99",X"B1",
		X"02",X"88",X"10",X"F7",X"4C",X"4D",X"EF",X"42",X"4C",X"4F",X"43",X"4B",X"53",X"20",X"46",X"52",
		X"45",X"45",X"2E",X"20",X"98",X"C3",X"20",X"20",X"C3",X"20",X"CA",X"C3",X"A9",X"00",X"85",X"86",
		X"20",X"9D",X"C4",X"30",X"3D",X"20",X"B7",X"DD",X"90",X"33",X"A0",X"00",X"B1",X"94",X"29",X"40",
		X"D0",X"2B",X"20",X"B6",X"C8",X"A0",X"13",X"B1",X"94",X"F0",X"0A",X"85",X"80",X"C8",X"B1",X"94",
		X"85",X"81",X"20",X"7D",X"C8",X"AE",X"53",X"02",X"A9",X"20",X"35",X"E7",X"D0",X"0D",X"BD",X"80",
		X"02",X"85",X"80",X"BD",X"85",X"02",X"85",X"81",X"20",X"7D",X"C8",X"E6",X"86",X"20",X"8B",X"C4",
		X"10",X"C3",X"A5",X"86",X"85",X"80",X"A9",X"01",X"A0",X"00",X"4C",X"A3",X"C1",X"20",X"5F",X"EF",
		X"20",X"75",X"D4",X"20",X"19",X"F1",X"B5",X"A7",X"C9",X"FF",X"F0",X"08",X"AD",X"F9",X"02",X"09",
		X"40",X"8D",X"F9",X"02",X"A9",X"00",X"20",X"C8",X"D4",X"20",X"56",X"D1",X"85",X"80",X"20",X"56",
		X"D1",X"85",X"81",X"A5",X"80",X"D0",X"06",X"20",X"F4",X"EE",X"4C",X"27",X"D2",X"20",X"5F",X"EF",
		X"20",X"4D",X"D4",X"4C",X"94",X"C8",X"A0",X"00",X"98",X"91",X"94",X"20",X"5E",X"DE",X"4C",X"99",
		X"D5",X"A9",X"31",X"4C",X"C8",X"C1",X"A9",X"4C",X"8D",X"00",X"06",X"A9",X"C7",X"8D",X"01",X"06",
		X"A9",X"FA",X"8D",X"02",X"06",X"A9",X"03",X"20",X"D3",X"D6",X"A5",X"7F",X"09",X"E0",X"85",X"03",
		X"A5",X"03",X"30",X"FC",X"C9",X"02",X"90",X"07",X"A9",X"03",X"A2",X"00",X"4C",X"0A",X"E6",X"60",
		X"A9",X"E0",X"8D",X"4F",X"02",X"20",X"D1",X"F0",X"20",X"19",X"F1",X"A9",X"FF",X"95",X"A7",X"A9",
		X"0F",X"8D",X"56",X"02",X"20",X"E5",X"C1",X"D0",X"03",X"4C",X"C1",X"C8",X"20",X"F8",X"C1",X"20",
		X"20",X"C3",X"AD",X"8B",X"02",X"29",X"55",X"D0",X"0F",X"AE",X"7A",X"02",X"BD",X"00",X"02",X"C9",
		X"2A",X"D0",X"05",X"A9",X"30",X"4C",X"C8",X"C1",X"AD",X"8B",X"02",X"29",X"D9",X"D0",X"F4",X"4C",
		X"52",X"C9",X"A9",X"00",X"8D",X"58",X"02",X"8D",X"8C",X"02",X"8D",X"80",X"02",X"8D",X"81",X"02",
		X"A5",X"E3",X"29",X"01",X"85",X"7F",X"09",X"01",X"8D",X"91",X"02",X"AD",X"7B",X"02",X"8D",X"7A",
		X"02",X"60",X"20",X"4F",X"C4",X"AD",X"78",X"02",X"C9",X"03",X"90",X"45",X"A5",X"E2",X"C5",X"E3",
		X"D0",X"3F",X"A5",X"DD",X"C5",X"DE",X"D0",X"39",X"A5",X"D8",X"C5",X"D9",X"D0",X"33",X"20",X"CC",
		X"CA",X"A9",X"01",X"8D",X"79",X"02",X"20",X"FA",X"C9",X"20",X"25",X"D1",X"F0",X"04",X"C9",X"02",
		X"D0",X"05",X"A9",X"64",X"20",X"C8",X"C1",X"A9",X"12",X"85",X"83",X"AD",X"3C",X"02",X"8D",X"3D",
		X"02",X"A9",X"FF",X"8D",X"3C",X"02",X"20",X"2A",X"DA",X"A2",X"02",X"20",X"B9",X"C9",X"4C",X"94",
		X"C1",X"20",X"A7",X"C9",X"4C",X"94",X"C1",X"20",X"E7",X"CA",X"A5",X"E2",X"29",X"01",X"85",X"7F",
		X"20",X"86",X"D4",X"20",X"E4",X"D6",X"AE",X"77",X"02",X"8E",X"79",X"02",X"20",X"FA",X"C9",X"A9",
		X"11",X"85",X"83",X"20",X"EB",X"D0",X"20",X"25",X"D1",X"D0",X"03",X"20",X"53",X"CA",X"A9",X"08",
		X"85",X"F8",X"4C",X"D8",X"C9",X"20",X"9B",X"CF",X"20",X"35",X"CA",X"A9",X"80",X"20",X"A6",X"DD",
		X"F0",X"F3",X"20",X"25",X"D1",X"F0",X"03",X"20",X"9B",X"CF",X"AE",X"79",X"02",X"E8",X"EC",X"78",
		X"02",X"90",X"C6",X"A9",X"12",X"85",X"83",X"4C",X"02",X"DB",X"AE",X"79",X"02",X"B5",X"E2",X"29",
		X"01",X"85",X"7F",X"AD",X"85",X"FE",X"85",X"80",X"B5",X"D8",X"85",X"81",X"20",X"75",X"D4",X"AE",
		X"79",X"02",X"B5",X"DD",X"20",X"C8",X"D4",X"AE",X"79",X"02",X"B5",X"E7",X"29",X"07",X"8D",X"4A",
		X"02",X"A9",X"00",X"8D",X"58",X"02",X"20",X"A0",X"D9",X"A0",X"01",X"20",X"25",X"D1",X"F0",X"01",
		X"C8",X"98",X"4C",X"C8",X"D4",X"A9",X"11",X"85",X"83",X"20",X"9B",X"D3",X"85",X"85",X"A6",X"82",
		X"B5",X"F2",X"29",X"08",X"85",X"F8",X"D0",X"0A",X"20",X"25",X"D1",X"F0",X"05",X"A9",X"80",X"20",
		X"97",X"DD",X"60",X"20",X"D3",X"D1",X"20",X"CB",X"E1",X"A5",X"D6",X"48",X"A5",X"D5",X"48",X"A9",
		X"12",X"85",X"83",X"20",X"07",X"D1",X"20",X"D3",X"D1",X"20",X"CB",X"E1",X"20",X"9C",X"E2",X"A5",
		X"D6",X"85",X"87",X"A5",X"D5",X"85",X"86",X"A9",X"00",X"85",X"88",X"85",X"D4",X"85",X"D7",X"68",
		X"85",X"D5",X"68",X"85",X"D6",X"4C",X"3B",X"E3",X"20",X"20",X"C3",X"A5",X"E3",X"29",X"01",X"85",
		X"E3",X"C5",X"E2",X"F0",X"02",X"09",X"80",X"85",X"E2",X"20",X"4F",X"C4",X"20",X"E7",X"CA",X"A5",
		X"E3",X"29",X"01",X"85",X"7F",X"A5",X"D9",X"85",X"81",X"20",X"57",X"DE",X"20",X"99",X"D5",X"A5",
		X"DE",X"18",X"69",X"03",X"20",X"C8",X"D4",X"20",X"93",X"DF",X"A8",X"AE",X"7A",X"02",X"A9",X"10",
		X"20",X"6E",X"C6",X"20",X"5E",X"DE",X"20",X"99",X"D5",X"4C",X"94",X"C1",X"A5",X"E8",X"29",X"07",
		X"8D",X"4A",X"02",X"AE",X"78",X"02",X"CA",X"EC",X"77",X"02",X"90",X"0A",X"BD",X"80",X"02",X"D0",
		X"F5",X"A9",X"62",X"4C",X"C8",X"C1",X"60",X"20",X"CC",X"CA",X"BD",X"80",X"02",X"F0",X"05",X"A9",
		X"63",X"4C",X"C8",X"C1",X"CA",X"10",X"F3",X"60",X"AD",X"01",X"02",X"C9",X"2D",X"D0",X"4C",X"AD",
		X"03",X"02",X"85",X"6F",X"AD",X"04",X"02",X"85",X"70",X"A0",X"00",X"AD",X"02",X"02",X"C9",X"52",
		X"F0",X"0E",X"20",X"58",X"F2",X"C9",X"57",X"F0",X"37",X"C9",X"45",X"D0",X"2E",X"6C",X"6F",X"00",
		X"B1",X"6F",X"85",X"85",X"AD",X"74",X"02",X"C9",X"06",X"90",X"1A",X"AE",X"05",X"02",X"CA",X"F0",
		X"14",X"8A",X"18",X"65",X"6F",X"E6",X"6F",X"8D",X"49",X"02",X"A5",X"6F",X"85",X"A5",X"A5",X"70",
		X"85",X"A6",X"4C",X"43",X"D4",X"20",X"EB",X"D0",X"4C",X"3A",X"D4",X"A9",X"31",X"4C",X"C8",X"C1",
		X"B9",X"06",X"02",X"91",X"6F",X"C8",X"CC",X"05",X"02",X"90",X"F5",X"60",X"AC",X"01",X"02",X"C0",
		X"30",X"D0",X"09",X"A9",X"EA",X"85",X"6B",X"A9",X"FF",X"85",X"6C",X"60",X"20",X"72",X"CB",X"4C",
		X"94",X"C1",X"88",X"98",X"29",X"0F",X"0A",X"A8",X"B1",X"6B",X"85",X"75",X"C8",X"B1",X"6B",X"85",
		X"76",X"6C",X"75",X"00",X"AD",X"8E",X"02",X"85",X"7F",X"A5",X"83",X"48",X"20",X"3D",X"C6",X"68",
		X"85",X"83",X"AE",X"74",X"02",X"CA",X"D0",X"0D",X"A9",X"01",X"20",X"E2",X"D1",X"4C",X"F1",X"CB",
		X"A9",X"70",X"4C",X"C8",X"C1",X"A0",X"01",X"20",X"7C",X"CC",X"AE",X"85",X"02",X"E0",X"05",X"B0",
		X"EF",X"A9",X"00",X"85",X"6F",X"85",X"70",X"38",X"26",X"6F",X"26",X"70",X"CA",X"10",X"F9",X"A5",
		X"6F",X"2D",X"4F",X"02",X"D0",X"DA",X"A5",X"70",X"2D",X"50",X"02",X"D0",X"D3",X"A5",X"6F",X"0D",
		X"4F",X"02",X"8D",X"4F",X"02",X"A5",X"70",X"0D",X"50",X"02",X"8D",X"50",X"02",X"A9",X"00",X"20",
		X"E2",X"D1",X"A6",X"82",X"AD",X"85",X"02",X"95",X"A7",X"AA",X"A5",X"7F",X"95",X"00",X"9D",X"5B",
		X"02",X"A6",X"83",X"BD",X"2B",X"02",X"09",X"40",X"9D",X"2B",X"02",X"A4",X"82",X"A9",X"FF",X"99",
		X"44",X"02",X"A9",X"89",X"99",X"F2",X"00",X"B9",X"A7",X"00",X"99",X"3E",X"02",X"0A",X"AA",X"A9",
		X"01",X"95",X"99",X"A9",X"0E",X"99",X"EC",X"00",X"4C",X"94",X"C1",X"A0",X"00",X"A2",X"00",X"A9",
		X"2D",X"20",X"68",X"C2",X"D0",X"0A",X"A9",X"31",X"4C",X"C8",X"C1",X"A9",X"30",X"4C",X"C8",X"C1",
		X"8A",X"D0",X"F8",X"A2",X"05",X"B9",X"00",X"02",X"DD",X"5D",X"CC",X"F0",X"05",X"CA",X"10",X"F8",
		X"30",X"E4",X"8A",X"09",X"80",X"8D",X"2A",X"02",X"20",X"6F",X"CC",X"AD",X"2A",X"02",X"0A",X"AA",
		X"BD",X"64",X"CC",X"85",X"70",X"BD",X"63",X"CC",X"85",X"6F",X"6C",X"6F",X"00",X"41",X"46",X"52",
		X"57",X"45",X"50",X"03",X"CD",X"F5",X"CC",X"56",X"CD",X"73",X"CD",X"A3",X"CD",X"BD",X"CD",X"A0",
		X"00",X"A2",X"00",X"A9",X"3A",X"20",X"68",X"C2",X"D0",X"02",X"A0",X"03",X"B9",X"00",X"02",X"C9",
		X"20",X"F0",X"08",X"C9",X"1D",X"F0",X"04",X"C9",X"2C",X"D0",X"07",X"C8",X"CC",X"74",X"02",X"90",
		X"EB",X"60",X"20",X"A1",X"CC",X"EE",X"77",X"02",X"AC",X"79",X"02",X"E0",X"04",X"90",X"EC",X"B0",
		X"8A",X"A9",X"00",X"85",X"6F",X"85",X"70",X"85",X"72",X"A2",X"FF",X"B9",X"00",X"02",X"C9",X"40",
		X"B0",X"18",X"C9",X"30",X"90",X"14",X"29",X"0F",X"48",X"A5",X"70",X"85",X"71",X"A5",X"6F",X"85",
		X"70",X"68",X"85",X"6F",X"C8",X"CC",X"74",X"02",X"90",X"E1",X"8C",X"79",X"02",X"18",X"A9",X"00",
		X"E8",X"E0",X"03",X"B0",X"0F",X"B4",X"6F",X"88",X"30",X"F6",X"7D",X"F2",X"CC",X"90",X"F8",X"18",
		X"E6",X"72",X"D0",X"F3",X"48",X"AE",X"77",X"02",X"A5",X"72",X"9D",X"80",X"02",X"68",X"9D",X"85",
		X"02",X"60",X"01",X"0A",X"64",X"20",X"F5",X"CD",X"20",X"5F",X"EF",X"4C",X"94",X"C1",X"A9",X"01",
		X"8D",X"F9",X"02",X"20",X"F5",X"CD",X"A5",X"81",X"48",X"20",X"FA",X"F1",X"F0",X"0B",X"68",X"C5",
		X"81",X"D0",X"19",X"20",X"90",X"EF",X"4C",X"94",X"C1",X"68",X"A9",X"00",X"85",X"81",X"E6",X"80",
		X"A5",X"80",X"CD",X"D7",X"FE",X"B0",X"0A",X"20",X"FA",X"F1",X"F0",X"EE",X"A9",X"65",X"20",X"45",
		X"E6",X"A9",X"65",X"20",X"C8",X"C1",X"20",X"F2",X"CD",X"4C",X"60",X"D4",X"20",X"2F",X"D1",X"A1",
		X"99",X"60",X"20",X"36",X"CD",X"A9",X"00",X"20",X"C8",X"D4",X"20",X"3C",X"CD",X"99",X"44",X"02",
		X"A9",X"89",X"99",X"F2",X"00",X"60",X"20",X"42",X"CD",X"20",X"EC",X"D3",X"4C",X"94",X"C1",X"20",
		X"6F",X"CC",X"20",X"42",X"CD",X"B9",X"44",X"02",X"99",X"3E",X"02",X"A9",X"FF",X"99",X"44",X"02",
		X"4C",X"94",X"C1",X"20",X"F2",X"CD",X"20",X"E8",X"D4",X"A8",X"88",X"C9",X"02",X"B0",X"02",X"A0",
		X"01",X"A9",X"00",X"20",X"C8",X"D4",X"98",X"20",X"F1",X"CF",X"8A",X"48",X"20",X"64",X"D4",X"68",
		X"AA",X"20",X"EE",X"D3",X"4C",X"94",X"C1",X"20",X"6F",X"CC",X"20",X"F2",X"CD",X"20",X"64",X"D4",
		X"4C",X"94",X"C1",X"20",X"58",X"F2",X"20",X"36",X"CD",X"A9",X"00",X"85",X"6F",X"A6",X"F9",X"BD",
		X"E0",X"FE",X"85",X"70",X"20",X"BA",X"CD",X"4C",X"94",X"C1",X"6C",X"6F",X"00",X"20",X"D2",X"CD",
		X"A5",X"F9",X"0A",X"AA",X"AD",X"86",X"02",X"95",X"99",X"20",X"2F",X"D1",X"20",X"EE",X"D3",X"4C",
		X"94",X"C1",X"A6",X"D3",X"E6",X"D3",X"BD",X"85",X"02",X"A8",X"88",X"88",X"C0",X"0C",X"90",X"05",
		X"A9",X"70",X"4C",X"C8",X"C1",X"85",X"83",X"20",X"EB",X"D0",X"B0",X"F4",X"20",X"93",X"DF",X"85",
		X"F9",X"60",X"20",X"D2",X"CD",X"A6",X"D3",X"BD",X"85",X"02",X"29",X"01",X"85",X"7F",X"BD",X"87",
		X"02",X"85",X"81",X"BD",X"86",X"02",X"85",X"80",X"20",X"5F",X"D5",X"4C",X"00",X"C1",X"20",X"2C",
		X"CE",X"20",X"6E",X"CE",X"A5",X"90",X"85",X"D7",X"20",X"71",X"CE",X"E6",X"D7",X"E6",X"D7",X"A5",
		X"8B",X"85",X"D5",X"A5",X"90",X"0A",X"18",X"69",X"10",X"85",X"D6",X"60",X"20",X"D9",X"CE",X"85",
		X"92",X"A6",X"82",X"B5",X"B5",X"85",X"90",X"B5",X"BB",X"85",X"91",X"D0",X"04",X"A5",X"90",X"F0",
		X"0B",X"A5",X"90",X"38",X"E9",X"01",X"85",X"90",X"B0",X"02",X"C6",X"91",X"B5",X"C7",X"85",X"6F",
		X"46",X"6F",X"90",X"03",X"20",X"ED",X"CE",X"20",X"E5",X"CE",X"A5",X"6F",X"D0",X"F2",X"A5",X"D4",
		X"18",X"65",X"8B",X"85",X"8B",X"90",X"06",X"E6",X"8C",X"D0",X"02",X"E6",X"8D",X"60",X"A9",X"FE",
		X"2C",X"A9",X"78",X"85",X"6F",X"A2",X"03",X"B5",X"8F",X"48",X"B5",X"8A",X"95",X"8F",X"68",X"95",
		X"8A",X"CA",X"D0",X"F3",X"20",X"D9",X"CE",X"A2",X"00",X"B5",X"90",X"95",X"8F",X"E8",X"E0",X"04",
		X"90",X"F7",X"A9",X"00",X"85",X"92",X"24",X"6F",X"30",X"09",X"06",X"8F",X"08",X"46",X"8F",X"28",
		X"20",X"E6",X"CE",X"20",X"ED",X"CE",X"20",X"E5",X"CE",X"24",X"6F",X"30",X"03",X"20",X"E2",X"CE",
		X"A5",X"8F",X"18",X"65",X"90",X"85",X"90",X"90",X"06",X"E6",X"91",X"D0",X"02",X"E6",X"92",X"A5",
		X"92",X"05",X"91",X"D0",X"C2",X"A5",X"90",X"38",X"E5",X"6F",X"90",X"0C",X"E6",X"8B",X"D0",X"06",
		X"E6",X"8C",X"D0",X"02",X"E6",X"8D",X"85",X"90",X"60",X"A9",X"00",X"85",X"8B",X"85",X"8C",X"85",
		X"8D",X"60",X"20",X"E5",X"CE",X"18",X"26",X"90",X"26",X"91",X"26",X"92",X"60",X"18",X"A2",X"FD",
		X"B5",X"8E",X"75",X"93",X"95",X"8E",X"E8",X"D0",X"F7",X"60",X"A2",X"00",X"8A",X"95",X"FA",X"E8",
		X"E0",X"04",X"D0",X"F8",X"A9",X"06",X"95",X"FA",X"60",X"A0",X"04",X"A6",X"82",X"B9",X"FA",X"00",
		X"96",X"FA",X"C5",X"82",X"F0",X"07",X"88",X"30",X"E1",X"AA",X"4C",X"0D",X"CF",X"60",X"20",X"09",
		X"CF",X"20",X"B7",X"DF",X"D0",X"46",X"20",X"D3",X"D1",X"20",X"8E",X"D2",X"30",X"48",X"20",X"C2",
		X"DF",X"A5",X"80",X"48",X"A5",X"81",X"48",X"A9",X"01",X"20",X"F6",X"D4",X"85",X"81",X"A9",X"00",
		X"20",X"F6",X"D4",X"85",X"80",X"F0",X"1F",X"20",X"25",X"D1",X"F0",X"0B",X"20",X"AB",X"DD",X"D0",
		X"06",X"20",X"8C",X"CF",X"4C",X"5D",X"CF",X"20",X"8C",X"CF",X"20",X"57",X"DE",X"68",X"85",X"81",
		X"68",X"85",X"80",X"4C",X"6F",X"CF",X"68",X"85",X"81",X"68",X"85",X"80",X"20",X"8C",X"CF",X"20",
		X"93",X"DF",X"AA",X"4C",X"99",X"D5",X"A9",X"70",X"4C",X"C8",X"C1",X"20",X"09",X"CF",X"20",X"B7",
		X"DF",X"D0",X"08",X"20",X"8E",X"D2",X"30",X"EE",X"20",X"C2",X"DF",X"60",X"A6",X"82",X"B5",X"A7",
		X"49",X"80",X"95",X"A7",X"B5",X"AE",X"49",X"80",X"95",X"AE",X"60",X"A2",X"12",X"86",X"83",X"20",
		X"07",X"D1",X"20",X"00",X"C1",X"20",X"25",X"D1",X"90",X"05",X"A9",X"20",X"20",X"9D",X"DD",X"A5",
		X"83",X"C9",X"0F",X"F0",X"23",X"D0",X"08",X"A5",X"84",X"29",X"8F",X"C9",X"0F",X"B0",X"19",X"20",
		X"25",X"D1",X"B0",X"05",X"A5",X"85",X"4C",X"9D",X"D1",X"D0",X"03",X"4C",X"AB",X"E0",X"A5",X"85",
		X"20",X"F1",X"CF",X"A4",X"82",X"4C",X"EE",X"D3",X"A9",X"04",X"85",X"82",X"20",X"E8",X"D4",X"C9",
		X"2A",X"F0",X"05",X"A5",X"85",X"20",X"F1",X"CF",X"A5",X"F8",X"F0",X"01",X"60",X"EE",X"55",X"02",
		X"60",X"48",X"20",X"93",X"DF",X"10",X"06",X"68",X"A9",X"61",X"4C",X"C8",X"C1",X"0A",X"AA",X"68",
		X"81",X"99",X"F6",X"99",X"60",X"20",X"D1",X"C1",X"20",X"42",X"D0",X"4C",X"94",X"C1",X"20",X"0F",
		X"F1",X"A8",X"B6",X"A7",X"E0",X"FF",X"D0",X"14",X"48",X"20",X"8E",X"D2",X"AA",X"10",X"05",X"A9",
		X"70",X"20",X"48",X"E6",X"68",X"A8",X"8A",X"09",X"80",X"99",X"A7",X"00",X"8A",X"29",X"0F",X"85",
		X"F9",X"A2",X"00",X"86",X"81",X"AE",X"85",X"FE",X"86",X"80",X"20",X"D3",X"D6",X"A9",X"B0",X"4C",
		X"8C",X"D5",X"20",X"D1",X"F0",X"20",X"13",X"D3",X"20",X"0E",X"D0",X"A6",X"7F",X"A9",X"00",X"9D",
		X"51",X"02",X"8A",X"0A",X"AA",X"A5",X"16",X"95",X"12",X"A5",X"17",X"95",X"13",X"20",X"86",X"D5",
		X"A5",X"F9",X"0A",X"AA",X"A9",X"02",X"95",X"99",X"A1",X"99",X"A6",X"7F",X"9D",X"01",X"01",X"A9",
		X"00",X"95",X"1C",X"95",X"FF",X"20",X"3A",X"EF",X"A0",X"04",X"A9",X"00",X"AA",X"18",X"71",X"6D",
		X"90",X"01",X"E8",X"C8",X"C8",X"C8",X"C8",X"C0",X"48",X"F0",X"F8",X"C0",X"90",X"D0",X"EE",X"48",
		X"8A",X"A6",X"7F",X"9D",X"FC",X"02",X"68",X"9D",X"FA",X"02",X"60",X"20",X"D0",X"D6",X"20",X"C3",
		X"D0",X"20",X"99",X"D5",X"20",X"37",X"D1",X"85",X"80",X"20",X"37",X"D1",X"85",X"81",X"60",X"20",
		X"9B",X"D0",X"A5",X"80",X"D0",X"01",X"60",X"20",X"1E",X"CF",X"20",X"D0",X"D6",X"20",X"C3",X"D0",
		X"4C",X"1E",X"CF",X"A9",X"80",X"D0",X"02",X"A9",X"90",X"8D",X"4D",X"02",X"20",X"93",X"DF",X"AA",
		X"20",X"06",X"D5",X"8A",X"48",X"0A",X"AA",X"A9",X"00",X"95",X"99",X"20",X"25",X"D1",X"C9",X"04",
		X"B0",X"06",X"F6",X"B5",X"D0",X"02",X"F6",X"BB",X"68",X"AA",X"60",X"A5",X"83",X"C9",X"13",X"90",
		X"02",X"29",X"0F",X"C9",X"0F",X"D0",X"02",X"A9",X"10",X"AA",X"38",X"BD",X"2B",X"02",X"30",X"06",
		X"29",X"0F",X"85",X"82",X"AA",X"18",X"60",X"A5",X"83",X"C9",X"13",X"90",X"02",X"29",X"0F",X"AA",
		X"BD",X"2B",X"02",X"A8",X"0A",X"90",X"0A",X"30",X"0A",X"98",X"29",X"0F",X"85",X"82",X"AA",X"18",
		X"60",X"30",X"F6",X"38",X"60",X"A6",X"82",X"B5",X"EC",X"4A",X"29",X"07",X"C9",X"04",X"60",X"20",
		X"93",X"DF",X"0A",X"AA",X"A4",X"82",X"60",X"20",X"2F",X"D1",X"B9",X"44",X"02",X"F0",X"12",X"A1",
		X"99",X"48",X"B5",X"99",X"D9",X"44",X"02",X"D0",X"04",X"A9",X"FF",X"95",X"99",X"68",X"F6",X"99",
		X"60",X"A1",X"99",X"F6",X"99",X"60",X"20",X"37",X"D1",X"D0",X"36",X"85",X"85",X"B9",X"44",X"02",
		X"F0",X"08",X"A9",X"80",X"99",X"F2",X"00",X"A5",X"85",X"60",X"20",X"1E",X"CF",X"A9",X"00",X"20",
		X"C8",X"D4",X"20",X"37",X"D1",X"C9",X"00",X"F0",X"19",X"85",X"80",X"20",X"37",X"D1",X"85",X"81",
		X"20",X"1E",X"CF",X"20",X"D3",X"D1",X"20",X"D0",X"D6",X"20",X"C3",X"D0",X"20",X"1E",X"CF",X"A5",
		X"85",X"60",X"20",X"37",X"D1",X"A4",X"82",X"99",X"44",X"02",X"A5",X"85",X"60",X"20",X"F1",X"CF",
		X"F0",X"01",X"60",X"20",X"D3",X"D1",X"20",X"1E",X"F1",X"A9",X"00",X"20",X"C8",X"D4",X"A5",X"80",
		X"20",X"F1",X"CF",X"A5",X"81",X"20",X"F1",X"CF",X"20",X"C7",X"D0",X"20",X"1E",X"CF",X"20",X"D0",
		X"D6",X"A9",X"02",X"4C",X"C8",X"D4",X"85",X"6F",X"20",X"E8",X"D4",X"18",X"65",X"6F",X"95",X"99",
		X"85",X"94",X"60",X"20",X"93",X"DF",X"AA",X"BD",X"5B",X"02",X"29",X"01",X"85",X"7F",X"60",X"38",
		X"B0",X"01",X"18",X"08",X"85",X"6F",X"20",X"27",X"D2",X"20",X"7F",X"D3",X"85",X"82",X"A6",X"83",
		X"28",X"90",X"02",X"09",X"80",X"9D",X"2B",X"02",X"29",X"3F",X"A8",X"A9",X"FF",X"99",X"A7",X"00",
		X"99",X"AE",X"00",X"99",X"CD",X"00",X"C6",X"6F",X"30",X"1C",X"20",X"8E",X"D2",X"10",X"08",X"20",
		X"5A",X"D2",X"A9",X"70",X"4C",X"C8",X"C1",X"99",X"A7",X"00",X"C6",X"6F",X"30",X"08",X"20",X"8E",
		X"D2",X"30",X"EC",X"99",X"AE",X"00",X"60",X"A5",X"83",X"C9",X"0F",X"D0",X"01",X"60",X"A6",X"83",
		X"BD",X"2B",X"02",X"C9",X"FF",X"F0",X"22",X"29",X"3F",X"85",X"82",X"A9",X"FF",X"9D",X"2B",X"02",
		X"A6",X"82",X"A9",X"00",X"95",X"F2",X"20",X"5A",X"D2",X"A6",X"82",X"A9",X"01",X"CA",X"30",X"03",
		X"0A",X"D0",X"FA",X"0D",X"56",X"02",X"8D",X"56",X"02",X"60",X"A6",X"82",X"B5",X"A7",X"C9",X"FF",
		X"F0",X"09",X"48",X"A9",X"FF",X"95",X"A7",X"68",X"20",X"F3",X"D2",X"A6",X"82",X"B5",X"AE",X"C9",
		X"FF",X"F0",X"09",X"48",X"A9",X"FF",X"95",X"AE",X"68",X"20",X"F3",X"D2",X"A6",X"82",X"B5",X"CD",
		X"C9",X"FF",X"F0",X"09",X"48",X"A9",X"FF",X"95",X"CD",X"68",X"20",X"F3",X"D2",X"60",X"98",X"48",
		X"A0",X"01",X"20",X"BA",X"D2",X"10",X"0C",X"88",X"20",X"BA",X"D2",X"10",X"06",X"20",X"39",X"D3",
		X"AA",X"30",X"13",X"B5",X"00",X"30",X"FC",X"A5",X"7F",X"95",X"00",X"9D",X"5B",X"02",X"8A",X"0A",
		X"A8",X"A9",X"02",X"99",X"99",X"00",X"68",X"A8",X"8A",X"60",X"A2",X"07",X"B9",X"4F",X"02",X"3D",
		X"E9",X"EF",X"F0",X"04",X"CA",X"10",X"F5",X"60",X"B9",X"4F",X"02",X"5D",X"E9",X"EF",X"99",X"4F",
		X"02",X"8A",X"88",X"30",X"03",X"18",X"69",X"08",X"AA",X"60",X"A6",X"82",X"B5",X"A7",X"30",X"09",
		X"8A",X"18",X"69",X"07",X"AA",X"B5",X"A7",X"10",X"F0",X"C9",X"FF",X"F0",X"EC",X"48",X"A9",X"FF",
		X"95",X"A7",X"68",X"29",X"0F",X"A8",X"C8",X"A2",X"10",X"6E",X"50",X"02",X"6E",X"4F",X"02",X"88",
		X"D0",X"01",X"18",X"CA",X"10",X"F3",X"60",X"A9",X"0E",X"85",X"83",X"20",X"27",X"D2",X"C6",X"83",
		X"D0",X"F9",X"60",X"A9",X"0E",X"85",X"83",X"A6",X"83",X"BD",X"2B",X"02",X"C9",X"FF",X"F0",X"14",
		X"29",X"3F",X"85",X"82",X"20",X"93",X"DF",X"AA",X"BD",X"5B",X"02",X"29",X"01",X"C5",X"7F",X"D0",
		X"03",X"20",X"27",X"D2",X"C6",X"83",X"10",X"DF",X"60",X"A5",X"6F",X"48",X"A0",X"00",X"B6",X"FA",
		X"B5",X"A7",X"10",X"04",X"C9",X"FF",X"D0",X"16",X"8A",X"18",X"69",X"07",X"AA",X"B5",X"A7",X"10",
		X"04",X"C9",X"FF",X"D0",X"09",X"C8",X"C0",X"05",X"90",X"E4",X"A2",X"FF",X"D0",X"1C",X"86",X"6F",
		X"29",X"3F",X"AA",X"B5",X"00",X"30",X"FC",X"C9",X"02",X"90",X"08",X"A6",X"6F",X"E0",X"07",X"90",
		X"D7",X"B0",X"E2",X"A4",X"6F",X"A9",X"FF",X"99",X"A7",X"00",X"68",X"85",X"6F",X"8A",X"60",X"A0",
		X"00",X"A9",X"01",X"2C",X"56",X"02",X"D0",X"09",X"C8",X"0A",X"D0",X"F7",X"A9",X"70",X"4C",X"C8",
		X"C1",X"49",X"FF",X"2D",X"56",X"02",X"8D",X"56",X"02",X"98",X"60",X"20",X"EB",X"D0",X"20",X"00",
		X"C1",X"20",X"AA",X"D3",X"A6",X"82",X"BD",X"3E",X"02",X"60",X"A6",X"82",X"20",X"25",X"D1",X"D0",
		X"03",X"4C",X"20",X"E1",X"A5",X"83",X"C9",X"0F",X"F0",X"5A",X"B5",X"F2",X"29",X"08",X"D0",X"13",
		X"20",X"25",X"D1",X"C9",X"07",X"D0",X"07",X"A9",X"89",X"95",X"F2",X"4C",X"DE",X"D3",X"A9",X"00",
		X"95",X"F2",X"60",X"A5",X"83",X"F0",X"32",X"20",X"25",X"D1",X"C9",X"04",X"90",X"22",X"20",X"2F",
		X"D1",X"B5",X"99",X"D9",X"44",X"02",X"D0",X"04",X"A9",X"00",X"95",X"99",X"F6",X"99",X"A1",X"99",
		X"99",X"3E",X"02",X"B5",X"99",X"D9",X"44",X"02",X"D0",X"05",X"A9",X"81",X"99",X"F2",X"00",X"60",
		X"20",X"56",X"D1",X"A6",X"82",X"9D",X"3E",X"02",X"60",X"AD",X"54",X"02",X"F0",X"F2",X"20",X"67",
		X"ED",X"4C",X"03",X"D4",X"20",X"E8",X"D4",X"C9",X"D4",X"D0",X"18",X"A5",X"95",X"C9",X"02",X"D0",
		X"12",X"A9",X"0D",X"85",X"85",X"20",X"23",X"C1",X"A9",X"00",X"20",X"C1",X"E6",X"C6",X"A5",X"A9",
		X"80",X"D0",X"12",X"20",X"37",X"D1",X"85",X"85",X"D0",X"09",X"A9",X"D4",X"20",X"C8",X"D4",X"A9",
		X"02",X"95",X"9A",X"A9",X"88",X"85",X"F7",X"A5",X"85",X"8D",X"43",X"02",X"60",X"20",X"93",X"DF",
		X"0A",X"AA",X"A9",X"00",X"95",X"99",X"A1",X"99",X"F0",X"05",X"D6",X"99",X"4C",X"56",X"D1",X"60",
		X"A9",X"80",X"D0",X"02",X"A9",X"90",X"05",X"7F",X"8D",X"4D",X"02",X"A5",X"F9",X"20",X"D3",X"D6",
		X"A6",X"F9",X"4C",X"93",X"D5",X"A9",X"01",X"8D",X"4A",X"02",X"A9",X"11",X"85",X"83",X"20",X"46",
		X"DC",X"A9",X"02",X"4C",X"C8",X"D4",X"A9",X"12",X"85",X"83",X"4C",X"DA",X"DC",X"20",X"3B",X"DE",
		X"A9",X"01",X"85",X"6F",X"A5",X"69",X"48",X"A9",X"03",X"85",X"69",X"20",X"2D",X"F1",X"68",X"85",
		X"69",X"A9",X"00",X"20",X"C8",X"D4",X"A5",X"80",X"20",X"F1",X"CF",X"A5",X"81",X"20",X"F1",X"CF",
		X"20",X"C7",X"D0",X"20",X"99",X"D5",X"A9",X"00",X"20",X"C8",X"D4",X"20",X"F1",X"CF",X"D0",X"FB",
		X"20",X"F1",X"CF",X"A9",X"FF",X"4C",X"F1",X"CF",X"85",X"6F",X"20",X"93",X"DF",X"0A",X"AA",X"B5",
		X"9A",X"85",X"95",X"A5",X"6F",X"95",X"99",X"85",X"94",X"60",X"A9",X"11",X"85",X"83",X"20",X"27",
		X"D2",X"A9",X"12",X"85",X"83",X"4C",X"27",X"D2",X"20",X"93",X"DF",X"0A",X"AA",X"B5",X"9A",X"85",
		X"95",X"B5",X"99",X"85",X"94",X"60",X"85",X"71",X"20",X"93",X"DF",X"AA",X"BD",X"E0",X"FE",X"85",
		X"72",X"A0",X"00",X"B1",X"71",X"60",X"BD",X"5B",X"02",X"29",X"01",X"0D",X"4D",X"02",X"48",X"86",
		X"F9",X"8A",X"0A",X"AA",X"B5",X"07",X"8D",X"4D",X"02",X"B5",X"06",X"F0",X"2D",X"CD",X"D7",X"FE",
		X"B0",X"28",X"AA",X"68",X"48",X"29",X"F0",X"C9",X"90",X"D0",X"4F",X"68",X"48",X"4A",X"B0",X"05",
		X"AD",X"01",X"01",X"90",X"03",X"AD",X"02",X"01",X"F0",X"05",X"CD",X"D5",X"FE",X"D0",X"33",X"8A",
		X"20",X"4B",X"F2",X"CD",X"4D",X"02",X"F0",X"02",X"B0",X"30",X"20",X"52",X"D5",X"A9",X"66",X"4C",
		X"45",X"E6",X"A5",X"F9",X"0A",X"AA",X"B5",X"06",X"85",X"80",X"B5",X"07",X"85",X"81",X"60",X"A5",
		X"80",X"F0",X"EA",X"CD",X"D7",X"FE",X"B0",X"E5",X"20",X"4B",X"F2",X"C5",X"81",X"F0",X"DE",X"90",
		X"DC",X"60",X"20",X"52",X"D5",X"A9",X"73",X"4C",X"45",X"E6",X"A6",X"F9",X"68",X"8D",X"4D",X"02",
		X"95",X"00",X"9D",X"5B",X"02",X"60",X"A9",X"80",X"D0",X"02",X"A9",X"90",X"05",X"7F",X"A6",X"F9",
		X"8D",X"4D",X"02",X"AD",X"4D",X"02",X"20",X"0E",X"D5",X"20",X"A6",X"D5",X"B0",X"FB",X"48",X"A9",
		X"00",X"8D",X"98",X"02",X"68",X"60",X"B5",X"00",X"30",X"1A",X"C9",X"02",X"90",X"14",X"C9",X"08",
		X"F0",X"08",X"C9",X"0B",X"F0",X"04",X"C9",X"0F",X"D0",X"0C",X"2C",X"98",X"02",X"30",X"03",X"4C",
		X"3F",X"D6",X"18",X"60",X"38",X"60",X"98",X"48",X"A5",X"7F",X"48",X"BD",X"5B",X"02",X"29",X"01",
		X"85",X"7F",X"A8",X"B9",X"CA",X"FE",X"8D",X"6D",X"02",X"20",X"A6",X"D6",X"C9",X"02",X"B0",X"03",
		X"4C",X"6D",X"D6",X"BD",X"5B",X"02",X"29",X"F0",X"48",X"C9",X"90",X"D0",X"07",X"A5",X"7F",X"09",
		X"B8",X"9D",X"5B",X"02",X"24",X"6A",X"70",X"39",X"A9",X"00",X"8D",X"99",X"02",X"8D",X"9A",X"02",
		X"AC",X"99",X"02",X"AD",X"9A",X"02",X"38",X"F9",X"DB",X"FE",X"8D",X"9A",X"02",X"B9",X"DB",X"FE",
		X"20",X"76",X"D6",X"EE",X"99",X"02",X"20",X"A6",X"D6",X"C9",X"02",X"90",X"08",X"AC",X"99",X"02",
		X"B9",X"DB",X"FE",X"D0",X"DB",X"AD",X"9A",X"02",X"20",X"76",X"D6",X"B5",X"00",X"C9",X"02",X"90",
		X"2B",X"24",X"6A",X"10",X"0F",X"68",X"C9",X"90",X"D0",X"05",X"05",X"7F",X"9D",X"5B",X"02",X"B5",
		X"00",X"20",X"0A",X"E6",X"68",X"2C",X"98",X"02",X"30",X"23",X"48",X"A9",X"C0",X"05",X"7F",X"95",
		X"00",X"B5",X"00",X"30",X"FC",X"20",X"A6",X"D6",X"C9",X"02",X"B0",X"D9",X"68",X"C9",X"90",X"D0",
		X"0C",X"05",X"7F",X"9D",X"5B",X"02",X"20",X"A6",X"D6",X"C9",X"02",X"B0",X"D2",X"68",X"85",X"7F",
		X"68",X"A8",X"B5",X"00",X"18",X"60",X"C9",X"00",X"F0",X"18",X"30",X"0C",X"A0",X"01",X"20",X"93",
		X"D6",X"38",X"E9",X"01",X"D0",X"F6",X"F0",X"0A",X"A0",X"FF",X"20",X"93",X"D6",X"18",X"69",X"01",
		X"D0",X"F6",X"60",X"48",X"98",X"A4",X"7F",X"99",X"FE",X"02",X"D9",X"FE",X"02",X"F0",X"FB",X"A9",
		X"00",X"99",X"FE",X"02",X"68",X"60",X"A5",X"6A",X"29",X"3F",X"A8",X"AD",X"6D",X"02",X"4D",X"00",
		X"1C",X"8D",X"00",X"1C",X"BD",X"5B",X"02",X"95",X"00",X"B5",X"00",X"30",X"FC",X"C9",X"02",X"90",
		X"03",X"88",X"D0",X"E7",X"48",X"AD",X"6D",X"02",X"0D",X"00",X"1C",X"8D",X"00",X"1C",X"68",X"60",
		X"20",X"93",X"DF",X"0A",X"A8",X"A5",X"80",X"99",X"06",X"00",X"A5",X"81",X"99",X"07",X"00",X"A5",
		X"7F",X"0A",X"AA",X"60",X"A5",X"83",X"48",X"A5",X"82",X"48",X"A5",X"81",X"48",X"A5",X"80",X"48",
		X"A9",X"11",X"85",X"83",X"20",X"3B",X"DE",X"AD",X"4A",X"02",X"48",X"A5",X"E2",X"29",X"01",X"85",
		X"7F",X"A6",X"F9",X"5D",X"5B",X"02",X"4A",X"90",X"0C",X"A2",X"01",X"8E",X"92",X"02",X"20",X"AC",
		X"C5",X"F0",X"1D",X"D0",X"28",X"AD",X"91",X"02",X"F0",X"0C",X"C5",X"81",X"F0",X"1F",X"85",X"81",
		X"20",X"60",X"D4",X"4C",X"3D",X"D7",X"A9",X"01",X"8D",X"92",X"02",X"20",X"17",X"C6",X"D0",X"0D",
		X"20",X"8D",X"D4",X"A5",X"81",X"8D",X"91",X"02",X"A9",X"02",X"8D",X"92",X"02",X"AD",X"92",X"02",
		X"20",X"C8",X"D4",X"68",X"8D",X"4A",X"02",X"C9",X"04",X"D0",X"02",X"09",X"80",X"20",X"F1",X"CF",
		X"68",X"8D",X"80",X"02",X"20",X"F1",X"CF",X"68",X"8D",X"85",X"02",X"20",X"F1",X"CF",X"20",X"93",
		X"DF",X"A8",X"AD",X"7A",X"02",X"AA",X"A9",X"10",X"20",X"6E",X"C6",X"A0",X"10",X"A9",X"00",X"91",
		X"94",X"C8",X"C0",X"1B",X"90",X"F9",X"AD",X"4A",X"02",X"C9",X"04",X"D0",X"13",X"A0",X"10",X"AD",
		X"59",X"02",X"91",X"94",X"C8",X"AD",X"5A",X"02",X"91",X"94",X"C8",X"AD",X"58",X"02",X"91",X"94",
		X"20",X"64",X"D4",X"68",X"85",X"82",X"AA",X"68",X"85",X"83",X"AD",X"91",X"02",X"85",X"D8",X"9D",
		X"60",X"02",X"AD",X"92",X"02",X"85",X"DD",X"9D",X"66",X"02",X"AD",X"4A",X"02",X"85",X"E7",X"A5",
		X"7F",X"85",X"E2",X"60",X"A5",X"83",X"8D",X"4C",X"02",X"20",X"B3",X"C2",X"8E",X"2A",X"02",X"AE",
		X"00",X"02",X"AD",X"4C",X"02",X"D0",X"2C",X"E0",X"2A",X"D0",X"28",X"A5",X"7E",X"F0",X"4D",X"85",
		X"80",X"AD",X"6E",X"02",X"85",X"7F",X"85",X"E2",X"A9",X"02",X"85",X"E7",X"AD",X"6F",X"02",X"85",
		X"81",X"20",X"00",X"C1",X"20",X"46",X"DC",X"A9",X"04",X"05",X"7F",X"A6",X"82",X"99",X"EC",X"00",
		X"4C",X"94",X"C1",X"E0",X"24",X"D0",X"1E",X"AD",X"4C",X"02",X"D0",X"03",X"4C",X"55",X"DA",X"20",
		X"D1",X"C1",X"AD",X"85",X"FE",X"85",X"80",X"A9",X"00",X"85",X"81",X"20",X"46",X"DC",X"A5",X"7F",
		X"09",X"02",X"4C",X"EB",X"D7",X"E0",X"23",X"D0",X"12",X"4C",X"84",X"CB",X"A9",X"02",X"8D",X"96",
		X"02",X"A9",X"00",X"85",X"7F",X"8D",X"8E",X"02",X"20",X"42",X"D0",X"20",X"E5",X"C1",X"D0",X"04",
		X"A2",X"00",X"F0",X"0C",X"8A",X"F0",X"05",X"A9",X"30",X"4C",X"C8",X"C1",X"88",X"F0",X"01",X"88",
		X"8C",X"7A",X"02",X"A9",X"8D",X"20",X"68",X"C2",X"E8",X"8E",X"78",X"02",X"20",X"12",X"C3",X"20",
		X"CA",X"C3",X"20",X"9D",X"C4",X"A2",X"00",X"8E",X"58",X"02",X"8E",X"97",X"02",X"8E",X"4A",X"02",
		X"E8",X"EC",X"77",X"02",X"B0",X"10",X"20",X"09",X"DA",X"E8",X"EC",X"77",X"02",X"B0",X"07",X"C0",
		X"04",X"F0",X"3E",X"20",X"09",X"DA",X"AE",X"4C",X"02",X"86",X"83",X"E0",X"02",X"B0",X"12",X"8E",
		X"97",X"02",X"A9",X"40",X"8D",X"F9",X"02",X"AD",X"4A",X"02",X"D0",X"1B",X"A9",X"02",X"8D",X"4A",
		X"02",X"AD",X"4A",X"02",X"D0",X"11",X"A5",X"E7",X"29",X"07",X"8D",X"4A",X"02",X"AD",X"80",X"02",
		X"D0",X"05",X"A9",X"01",X"8D",X"4A",X"02",X"AD",X"97",X"02",X"C9",X"01",X"F0",X"18",X"4C",X"40",
		X"D9",X"BC",X"7A",X"02",X"B9",X"00",X"02",X"8D",X"58",X"02",X"AD",X"80",X"02",X"D0",X"B7",X"A9",
		X"01",X"8D",X"97",X"02",X"D0",X"B0",X"A5",X"E7",X"29",X"80",X"AA",X"D0",X"14",X"A9",X"20",X"24",
		X"E7",X"F0",X"06",X"20",X"B6",X"C8",X"4C",X"E3",X"D9",X"AD",X"80",X"02",X"D0",X"03",X"4C",X"E3",
		X"D9",X"AD",X"00",X"02",X"C9",X"40",X"F0",X"0D",X"8A",X"D0",X"05",X"A9",X"63",X"4C",X"C8",X"C1",
		X"A9",X"33",X"4C",X"C8",X"C1",X"A5",X"E7",X"29",X"07",X"CD",X"4A",X"02",X"D0",X"67",X"C9",X"04",
		X"F0",X"63",X"20",X"DA",X"DC",X"A5",X"82",X"8D",X"70",X"02",X"A9",X"11",X"85",X"83",X"20",X"EB",
		X"D0",X"AD",X"94",X"02",X"20",X"C8",X"D4",X"A0",X"00",X"B1",X"94",X"09",X"20",X"91",X"94",X"A0",
		X"1A",X"A5",X"80",X"91",X"94",X"C8",X"A5",X"81",X"91",X"94",X"AE",X"70",X"02",X"A5",X"D8",X"9D",
		X"60",X"02",X"A5",X"DD",X"9D",X"66",X"02",X"20",X"3B",X"DE",X"20",X"64",X"D4",X"4C",X"EF",X"D9",
		X"AD",X"80",X"02",X"D0",X"05",X"A9",X"62",X"4C",X"C8",X"C1",X"AD",X"97",X"02",X"C9",X"03",X"F0",
		X"0B",X"A9",X"20",X"24",X"E7",X"F0",X"05",X"A9",X"60",X"4C",X"C8",X"C1",X"A5",X"E7",X"29",X"07",
		X"CD",X"4A",X"02",X"F0",X"05",X"A9",X"64",X"4C",X"C8",X"C1",X"A0",X"00",X"8C",X"79",X"02",X"AE",
		X"97",X"02",X"E0",X"02",X"D0",X"1A",X"C9",X"04",X"F0",X"EB",X"B1",X"94",X"29",X"4F",X"91",X"94",
		X"A5",X"83",X"48",X"A9",X"11",X"85",X"83",X"20",X"3B",X"DE",X"20",X"64",X"D4",X"68",X"85",X"83",
		X"20",X"A0",X"D9",X"AD",X"97",X"02",X"C9",X"02",X"D0",X"55",X"20",X"2A",X"DA",X"4C",X"94",X"C1",
		X"A0",X"13",X"B1",X"94",X"8D",X"59",X"02",X"C8",X"B1",X"94",X"8D",X"5A",X"02",X"C8",X"B1",X"94",
		X"AE",X"58",X"02",X"8D",X"58",X"02",X"8A",X"F0",X"0A",X"CD",X"58",X"02",X"F0",X"05",X"A9",X"50",
		X"20",X"C8",X"C1",X"AE",X"79",X"02",X"BD",X"80",X"02",X"85",X"80",X"BD",X"85",X"02",X"85",X"81",
		X"20",X"46",X"DC",X"A4",X"82",X"AE",X"79",X"02",X"B5",X"D8",X"99",X"60",X"02",X"B5",X"DD",X"99",
		X"66",X"02",X"60",X"A5",X"E2",X"29",X"01",X"85",X"7F",X"20",X"DA",X"DC",X"20",X"E4",X"D6",X"A5",
		X"83",X"C9",X"02",X"B0",X"11",X"20",X"3E",X"DE",X"A5",X"80",X"85",X"7E",X"A5",X"7F",X"8D",X"6E",
		X"02",X"A5",X"81",X"8D",X"6F",X"02",X"4C",X"99",X"C1",X"BC",X"7A",X"02",X"B9",X"00",X"02",X"A0",
		X"04",X"88",X"30",X"08",X"D9",X"B2",X"FE",X"D0",X"F8",X"8C",X"97",X"02",X"A0",X"05",X"88",X"30",
		X"08",X"D9",X"B6",X"FE",X"D0",X"F8",X"8C",X"4A",X"02",X"60",X"20",X"39",X"CA",X"A9",X"80",X"20",
		X"A6",X"DD",X"F0",X"F6",X"20",X"95",X"DE",X"A6",X"81",X"E8",X"8A",X"D0",X"05",X"20",X"A3",X"D1",
		X"A9",X"02",X"20",X"C8",X"D4",X"A6",X"82",X"A9",X"01",X"95",X"F2",X"A9",X"80",X"05",X"82",X"A6",
		X"83",X"9D",X"2B",X"02",X"60",X"A9",X"0C",X"8D",X"2A",X"02",X"A9",X"00",X"AE",X"74",X"02",X"CA",
		X"F0",X"0B",X"CA",X"D0",X"21",X"AD",X"01",X"02",X"20",X"BD",X"C3",X"30",X"19",X"85",X"E2",X"EE",
		X"77",X"02",X"EE",X"78",X"02",X"EE",X"7A",X"02",X"A9",X"80",X"85",X"E7",X"A9",X"2A",X"8D",X"00",
		X"02",X"8D",X"01",X"02",X"D0",X"18",X"20",X"E5",X"C1",X"D0",X"05",X"20",X"DC",X"C2",X"A0",X"03",
		X"88",X"88",X"8C",X"7A",X"02",X"20",X"00",X"C2",X"20",X"98",X"C3",X"20",X"20",X"C3",X"20",X"CA",
		X"C3",X"20",X"B7",X"C7",X"20",X"9D",X"C4",X"20",X"9E",X"EC",X"20",X"37",X"D1",X"A6",X"82",X"9D",
		X"3E",X"02",X"A5",X"7F",X"8D",X"8E",X"02",X"09",X"04",X"95",X"EC",X"A9",X"00",X"85",X"A3",X"60",
		X"A9",X"00",X"8D",X"F9",X"02",X"A5",X"83",X"D0",X"0B",X"A9",X"00",X"8D",X"54",X"02",X"20",X"27",
		X"D2",X"4C",X"DA",X"D4",X"C9",X"0F",X"F0",X"14",X"20",X"02",X"DB",X"A5",X"83",X"C9",X"02",X"90",
		X"F0",X"AD",X"6C",X"02",X"D0",X"03",X"4C",X"94",X"C1",X"4C",X"AD",X"C1",X"A9",X"0E",X"85",X"83",
		X"20",X"02",X"DB",X"C6",X"83",X"10",X"F9",X"AD",X"6C",X"02",X"D0",X"03",X"4C",X"94",X"C1",X"4C",
		X"AD",X"C1",X"A6",X"83",X"BD",X"2B",X"02",X"C9",X"FF",X"D0",X"01",X"60",X"29",X"0F",X"85",X"82",
		X"20",X"25",X"D1",X"C9",X"07",X"F0",X"0F",X"C9",X"04",X"F0",X"11",X"20",X"07",X"D1",X"B0",X"09",
		X"20",X"62",X"DB",X"20",X"A5",X"DB",X"20",X"F4",X"EE",X"4C",X"27",X"D2",X"20",X"F1",X"DD",X"20",
		X"1E",X"CF",X"20",X"CB",X"E1",X"A6",X"D5",X"86",X"73",X"E6",X"73",X"A9",X"00",X"85",X"70",X"85",
		X"71",X"A5",X"D6",X"38",X"E9",X"0E",X"85",X"72",X"20",X"51",X"DF",X"A6",X"82",X"A5",X"70",X"95",
		X"B5",X"A5",X"71",X"95",X"BB",X"A9",X"40",X"20",X"A6",X"DD",X"F0",X"03",X"20",X"A5",X"DB",X"4C",
		X"27",X"D2",X"A6",X"82",X"B5",X"B5",X"15",X"BB",X"D0",X"0C",X"20",X"E8",X"D4",X"C9",X"02",X"D0",
		X"05",X"A9",X"0D",X"20",X"F1",X"CF",X"20",X"E8",X"D4",X"C9",X"02",X"D0",X"0F",X"20",X"1E",X"CF",
		X"A6",X"82",X"B5",X"B5",X"D0",X"02",X"D6",X"BB",X"D6",X"B5",X"A9",X"00",X"38",X"E9",X"01",X"48",
		X"A9",X"00",X"20",X"C8",X"D4",X"20",X"F1",X"CF",X"68",X"20",X"F1",X"CF",X"20",X"C7",X"D0",X"20",
		X"99",X"D5",X"4C",X"1E",X"CF",X"A6",X"82",X"8E",X"70",X"02",X"A5",X"83",X"48",X"BD",X"60",X"02",
		X"85",X"81",X"BD",X"66",X"02",X"8D",X"94",X"02",X"B5",X"EC",X"29",X"01",X"85",X"7F",X"AD",X"85",
		X"FE",X"85",X"80",X"20",X"93",X"DF",X"48",X"85",X"F9",X"20",X"60",X"D4",X"A0",X"00",X"BD",X"E0",
		X"FE",X"85",X"87",X"AD",X"94",X"02",X"85",X"86",X"B1",X"86",X"29",X"20",X"F0",X"43",X"20",X"25",
		X"D1",X"C9",X"04",X"F0",X"44",X"B1",X"86",X"29",X"8F",X"91",X"86",X"C8",X"B1",X"86",X"85",X"80",
		X"84",X"71",X"A0",X"1B",X"B1",X"86",X"48",X"88",X"B1",X"86",X"D0",X"0A",X"85",X"80",X"68",X"85",
		X"81",X"A9",X"67",X"20",X"45",X"E6",X"48",X"A9",X"00",X"91",X"86",X"C8",X"91",X"86",X"68",X"A4",
		X"71",X"91",X"86",X"C8",X"B1",X"86",X"85",X"81",X"68",X"91",X"86",X"20",X"7D",X"C8",X"4C",X"29",
		X"DC",X"B1",X"86",X"29",X"0F",X"09",X"80",X"91",X"86",X"AE",X"70",X"02",X"A0",X"1C",X"B5",X"B5",
		X"91",X"86",X"C8",X"B5",X"BB",X"91",X"86",X"68",X"AA",X"A9",X"90",X"05",X"7F",X"20",X"90",X"D5",
		X"68",X"85",X"83",X"4C",X"07",X"D1",X"A9",X"01",X"20",X"E2",X"D1",X"20",X"B6",X"DC",X"AD",X"4A",
		X"02",X"48",X"0A",X"05",X"7F",X"95",X"EC",X"20",X"9B",X"D0",X"A6",X"82",X"A5",X"80",X"D0",X"05",
		X"A5",X"81",X"9D",X"44",X"02",X"68",X"C9",X"04",X"D0",X"3F",X"A4",X"83",X"B9",X"2B",X"02",X"09",
		X"40",X"99",X"2B",X"02",X"AD",X"58",X"02",X"95",X"C7",X"20",X"8E",X"D2",X"10",X"03",X"4C",X"0F",
		X"D2",X"A6",X"82",X"95",X"CD",X"AC",X"59",X"02",X"84",X"80",X"AC",X"5A",X"02",X"84",X"81",X"20",
		X"D3",X"D6",X"20",X"73",X"DE",X"20",X"99",X"D5",X"A6",X"82",X"A9",X"02",X"95",X"C1",X"A9",X"00",
		X"20",X"C8",X"D4",X"20",X"53",X"E1",X"4C",X"3E",X"DE",X"20",X"56",X"D1",X"A6",X"82",X"9D",X"3E",
		X"02",X"A9",X"88",X"95",X"F2",X"60",X"A6",X"82",X"B5",X"A7",X"0A",X"A8",X"A9",X"02",X"99",X"99",
		X"00",X"B5",X"AE",X"09",X"80",X"95",X"AE",X"0A",X"A8",X"A9",X"02",X"99",X"99",X"00",X"A9",X"00",
		X"95",X"B5",X"95",X"BB",X"A9",X"00",X"9D",X"44",X"02",X"60",X"20",X"A9",X"F1",X"A9",X"01",X"20",
		X"DF",X"D1",X"20",X"D0",X"D6",X"20",X"B6",X"DC",X"A6",X"82",X"AD",X"4A",X"02",X"48",X"0A",X"05",
		X"7F",X"95",X"EC",X"68",X"C9",X"04",X"F0",X"05",X"A9",X"01",X"95",X"F2",X"60",X"A4",X"83",X"B9",
		X"2B",X"02",X"29",X"3F",X"09",X"40",X"99",X"2B",X"02",X"AD",X"58",X"02",X"95",X"C7",X"20",X"8E",
		X"D2",X"10",X"03",X"4C",X"0F",X"D2",X"A6",X"82",X"95",X"CD",X"20",X"C1",X"DE",X"20",X"1E",X"F1",
		X"A5",X"80",X"8D",X"59",X"02",X"A5",X"81",X"8D",X"5A",X"02",X"A6",X"82",X"B5",X"CD",X"20",X"D3",
		X"D6",X"A9",X"00",X"20",X"E9",X"DE",X"A9",X"00",X"20",X"8D",X"DD",X"A9",X"11",X"20",X"8D",X"DD",
		X"A9",X"00",X"20",X"8D",X"DD",X"AD",X"58",X"02",X"20",X"8D",X"DD",X"A5",X"80",X"20",X"8D",X"DD",
		X"A5",X"81",X"20",X"8D",X"DD",X"A9",X"10",X"20",X"E9",X"DE",X"20",X"3E",X"DE",X"A5",X"80",X"20",
		X"8D",X"DD",X"A5",X"81",X"20",X"8D",X"DD",X"20",X"6C",X"DE",X"20",X"99",X"D5",X"A9",X"02",X"20",
		X"C8",X"D4",X"A6",X"82",X"38",X"A9",X"00",X"F5",X"C7",X"95",X"C1",X"20",X"E2",X"E2",X"20",X"19",
		X"DE",X"20",X"5E",X"DE",X"20",X"99",X"D5",X"20",X"F4",X"EE",X"4C",X"98",X"DC",X"48",X"A6",X"82",
		X"B5",X"CD",X"4C",X"FD",X"CF",X"90",X"06",X"A6",X"82",X"15",X"EC",X"D0",X"06",X"A6",X"82",X"49",
		X"FF",X"35",X"EC",X"95",X"EC",X"60",X"A6",X"82",X"35",X"EC",X"60",X"20",X"93",X"DF",X"AA",X"BD",
		X"5B",X"02",X"29",X"F0",X"C9",X"90",X"60",X"A2",X"00",X"86",X"71",X"BD",X"2B",X"02",X"C9",X"FF",
		X"D0",X"08",X"A6",X"71",X"E8",X"E0",X"10",X"90",X"F0",X"60",X"86",X"71",X"29",X"3F",X"A8",X"B9",
		X"EC",X"00",X"29",X"01",X"85",X"70",X"AE",X"53",X"02",X"B5",X"E2",X"29",X"01",X"C5",X"70",X"D0",
		X"E1",X"B9",X"60",X"02",X"D5",X"D8",X"D0",X"DA",X"B9",X"66",X"02",X"D5",X"DD",X"D0",X"D3",X"18",
		X"60",X"20",X"9E",X"DF",X"50",X"06",X"20",X"5E",X"DE",X"20",X"99",X"D5",X"60",X"20",X"2B",X"DE",
		X"A5",X"80",X"91",X"94",X"C8",X"A5",X"81",X"91",X"94",X"4C",X"05",X"E1",X"20",X"2B",X"DE",X"B1",
		X"94",X"85",X"80",X"C8",X"B1",X"94",X"85",X"81",X"60",X"20",X"2B",X"DE",X"A9",X"00",X"91",X"94",
		X"C8",X"A6",X"82",X"B5",X"C1",X"AA",X"CA",X"8A",X"91",X"94",X"60",X"20",X"93",X"DF",X"0A",X"AA",
		X"B5",X"9A",X"85",X"95",X"A9",X"00",X"85",X"94",X"A0",X"00",X"60",X"20",X"EB",X"D0",X"20",X"93",
		X"DF",X"85",X"F9",X"0A",X"A8",X"B9",X"06",X"00",X"85",X"80",X"B9",X"07",X"00",X"85",X"81",X"60",
		X"A9",X"90",X"8D",X"4D",X"02",X"D0",X"28",X"A9",X"80",X"8D",X"4D",X"02",X"D0",X"21",X"A9",X"90",
		X"8D",X"4D",X"02",X"D0",X"26",X"A9",X"80",X"8D",X"4D",X"02",X"D0",X"1F",X"A9",X"90",X"8D",X"4D",
		X"02",X"D0",X"02",X"A9",X"80",X"8D",X"4D",X"02",X"A6",X"82",X"B5",X"CD",X"AA",X"10",X"13",X"20",
		X"D0",X"D6",X"20",X"93",X"DF",X"AA",X"A5",X"7F",X"9D",X"5B",X"02",X"20",X"15",X"E1",X"20",X"93",
		X"DF",X"AA",X"4C",X"06",X"D5",X"A9",X"00",X"20",X"C8",X"D4",X"20",X"37",X"D1",X"85",X"80",X"20",
		X"37",X"D1",X"85",X"81",X"60",X"48",X"A9",X"00",X"85",X"6F",X"85",X"71",X"B9",X"E0",X"FE",X"85",
		X"70",X"BD",X"E0",X"FE",X"85",X"72",X"68",X"A8",X"88",X"B1",X"6F",X"91",X"71",X"88",X"10",X"F9",
		X"60",X"A8",X"B9",X"E0",X"FE",X"85",X"70",X"A9",X"00",X"85",X"6F",X"A8",X"91",X"6F",X"C8",X"D0",
		X"FB",X"60",X"A9",X"00",X"20",X"DC",X"DE",X"A0",X"02",X"B1",X"94",X"60",X"85",X"94",X"A6",X"82",
		X"B5",X"CD",X"AA",X"BD",X"E0",X"FE",X"85",X"95",X"60",X"48",X"20",X"DC",X"DE",X"48",X"8A",X"0A",
		X"AA",X"68",X"95",X"9A",X"68",X"95",X"99",X"60",X"20",X"66",X"DF",X"30",X"0E",X"50",X"13",X"A6",
		X"82",X"B5",X"CD",X"20",X"1B",X"DF",X"20",X"66",X"DF",X"10",X"07",X"20",X"CB",X"E1",X"2C",X"CE",
		X"FE",X"60",X"A5",X"D6",X"20",X"E9",X"DE",X"2C",X"CD",X"FE",X"60",X"85",X"F9",X"A9",X"80",X"D0",
		X"04",X"85",X"F9",X"A9",X"90",X"48",X"B5",X"EC",X"29",X"01",X"85",X"7F",X"68",X"05",X"7F",X"8D",
		X"4D",X"02",X"B1",X"94",X"85",X"80",X"C8",X"B1",X"94",X"85",X"81",X"A5",X"F9",X"20",X"D3",X"D6",
		X"A6",X"F9",X"4C",X"93",X"D5",X"A6",X"82",X"B5",X"CD",X"4C",X"EB",X"D4",X"A9",X"78",X"20",X"5C",
		X"DF",X"CA",X"10",X"F8",X"A5",X"72",X"4A",X"20",X"5C",X"DF",X"A5",X"73",X"18",X"65",X"70",X"85",
		X"70",X"90",X"02",X"E6",X"71",X"60",X"20",X"D2",X"DE",X"C5",X"D5",X"D0",X"0E",X"A4",X"D6",X"B1",
		X"94",X"F0",X"04",X"2C",X"CD",X"FE",X"60",X"2C",X"CF",X"FE",X"60",X"A5",X"D5",X"C9",X"06",X"B0",
		X"0A",X"0A",X"A8",X"A9",X"04",X"85",X"94",X"B1",X"94",X"D0",X"04",X"2C",X"D0",X"FE",X"60",X"2C",
		X"CE",X"FE",X"60",X"A6",X"82",X"B5",X"A7",X"10",X"02",X"B5",X"AE",X"29",X"BF",X"60",X"A6",X"82",
		X"8E",X"57",X"02",X"B5",X"A7",X"10",X"09",X"8A",X"18",X"69",X"07",X"8D",X"57",X"02",X"B5",X"AE",
		X"85",X"70",X"29",X"1F",X"24",X"70",X"60",X"A6",X"82",X"B5",X"A7",X"30",X"02",X"B5",X"AE",X"C9",
		X"FF",X"60",X"A6",X"82",X"09",X"80",X"B4",X"A7",X"10",X"03",X"95",X"A7",X"60",X"95",X"AE",X"60",
		X"A9",X"20",X"20",X"9D",X"DD",X"A9",X"80",X"20",X"A6",X"DD",X"D0",X"41",X"A6",X"82",X"F6",X"B5",
		X"D0",X"02",X"F6",X"BB",X"A6",X"82",X"B5",X"C1",X"F0",X"2E",X"20",X"E8",X"D4",X"A6",X"82",X"D5",
		X"C1",X"90",X"03",X"20",X"3C",X"E0",X"A6",X"82",X"B5",X"C1",X"20",X"C8",X"D4",X"A1",X"99",X"85",
		X"85",X"A9",X"20",X"20",X"9D",X"DD",X"20",X"04",X"E3",X"48",X"90",X"28",X"A9",X"00",X"20",X"F6",
		X"D4",X"D0",X"21",X"68",X"C9",X"02",X"F0",X"12",X"A9",X"80",X"20",X"97",X"DD",X"20",X"2F",X"D1",
		X"B5",X"99",X"99",X"44",X"02",X"A9",X"0D",X"85",X"85",X"60",X"20",X"35",X"E0",X"A6",X"82",X"A9",
		X"00",X"95",X"C1",X"60",X"68",X"A6",X"82",X"95",X"C1",X"4C",X"6E",X"E1",X"20",X"D3",X"D1",X"20",
		X"95",X"DE",X"20",X"9E",X"DF",X"50",X"16",X"20",X"5E",X"DE",X"20",X"1E",X"CF",X"A9",X"02",X"20",
		X"C8",X"D4",X"20",X"AB",X"DD",X"D0",X"24",X"20",X"57",X"DE",X"4C",X"99",X"D5",X"20",X"1E",X"CF",
		X"20",X"AB",X"DD",X"D0",X"06",X"20",X"57",X"DE",X"20",X"99",X"D5",X"20",X"95",X"DE",X"A5",X"80",
		X"F0",X"09",X"20",X"1E",X"CF",X"20",X"57",X"DE",X"20",X"1E",X"CF",X"60",X"20",X"05",X"E1",X"20",
		X"93",X"DF",X"0A",X"AA",X"A5",X"85",X"81",X"99",X"B4",X"99",X"C8",X"D0",X"09",X"A4",X"82",X"B9",
		X"C1",X"00",X"F0",X"0A",X"A0",X"02",X"98",X"A4",X"82",X"D9",X"C1",X"00",X"D0",X"05",X"A9",X"20",
		X"4C",X"97",X"DD",X"F6",X"99",X"D0",X"03",X"20",X"3C",X"E0",X"60",X"A9",X"A0",X"20",X"A6",X"DD",
		X"D0",X"27",X"A5",X"85",X"20",X"7C",X"E0",X"A5",X"F8",X"F0",X"0D",X"60",X"A9",X"20",X"20",X"A6",
		X"DD",X"F0",X"05",X"A9",X"51",X"8D",X"6C",X"02",X"20",X"F3",X"E0",X"20",X"53",X"E1",X"AD",X"6C",
		X"02",X"F0",X"03",X"4C",X"C8",X"C1",X"4C",X"BC",X"E6",X"29",X"80",X"D0",X"05",X"A5",X"F8",X"F0",
		X"DB",X"60",X"A5",X"85",X"48",X"20",X"1C",X"E3",X"68",X"85",X"85",X"A9",X"80",X"20",X"9D",X"DD",
		X"4C",X"B2",X"E0",X"A9",X"20",X"20",X"A6",X"DD",X"D0",X"0A",X"A9",X"00",X"85",X"85",X"20",X"7C",
		X"E0",X"4C",X"F3",X"E0",X"60",X"A9",X"40",X"20",X"97",X"DD",X"20",X"9E",X"DF",X"09",X"40",X"AE",
		X"57",X"02",X"95",X"A7",X"60",X"20",X"9E",X"DF",X"29",X"BF",X"AE",X"57",X"02",X"95",X"A7",X"60",
		X"A9",X"80",X"20",X"A6",X"DD",X"D0",X"37",X"20",X"2F",X"D1",X"B5",X"99",X"D9",X"44",X"02",X"F0",
		X"22",X"F6",X"99",X"D0",X"06",X"20",X"3C",X"E0",X"20",X"2F",X"D1",X"A1",X"99",X"99",X"3E",X"02",
		X"A9",X"89",X"99",X"F2",X"00",X"B5",X"99",X"D9",X"44",X"02",X"F0",X"01",X"60",X"A9",X"81",X"99",
		X"F2",X"00",X"60",X"20",X"D0",X"DF",X"20",X"2F",X"D1",X"A5",X"85",X"4C",X"3D",X"E1",X"A6",X"82",
		X"A9",X"0D",X"9D",X"3E",X"02",X"A9",X"81",X"95",X"F2",X"A9",X"50",X"20",X"C8",X"C1",X"A6",X"82",
		X"B5",X"C1",X"85",X"87",X"C6",X"87",X"C9",X"02",X"D0",X"04",X"A9",X"FF",X"85",X"87",X"B5",X"C7",
		X"85",X"88",X"20",X"E8",X"D4",X"A6",X"82",X"C5",X"87",X"90",X"19",X"F0",X"17",X"20",X"1E",X"CF",
		X"20",X"B2",X"E1",X"90",X"08",X"A6",X"82",X"9D",X"44",X"02",X"4C",X"1E",X"CF",X"20",X"1E",X"CF",
		X"A9",X"FF",X"85",X"87",X"20",X"B2",X"E1",X"B0",X"03",X"20",X"E8",X"D4",X"A6",X"82",X"9D",X"44",
		X"02",X"60",X"20",X"2B",X"DE",X"A4",X"87",X"B1",X"94",X"D0",X"0D",X"88",X"C0",X"02",X"90",X"04",
		X"C6",X"88",X"D0",X"F3",X"C6",X"88",X"18",X"60",X"98",X"38",X"60",X"20",X"D2",X"DE",X"85",X"D5",
		X"A9",X"04",X"85",X"94",X"A0",X"0A",X"D0",X"04",X"88",X"88",X"30",X"26",X"B1",X"94",X"F0",X"F8",
		X"98",X"4A",X"C5",X"D5",X"F0",X"09",X"85",X"D5",X"A6",X"82",X"B5",X"CD",X"20",X"1B",X"DF",X"A0",
		X"00",X"84",X"94",X"B1",X"94",X"D0",X"0B",X"C8",X"B1",X"94",X"A8",X"88",X"84",X"D6",X"98",X"4C",
		X"E9",X"DE",X"A9",X"67",X"20",X"45",X"E6",X"20",X"B3",X"C2",X"AD",X"01",X"02",X"85",X"83",X"20",
		X"EB",X"D0",X"90",X"05",X"A9",X"70",X"20",X"C8",X"C1",X"A9",X"A0",X"20",X"9D",X"DD",X"20",X"25",
		X"D1",X"F0",X"05",X"A9",X"64",X"20",X"C8",X"C1",X"B5",X"EC",X"29",X"01",X"85",X"7F",X"AD",X"02",
		X"02",X"95",X"B5",X"AD",X"03",X"02",X"95",X"BB",X"A6",X"82",X"A9",X"89",X"95",X"F2",X"AD",X"04",
		X"02",X"F0",X"10",X"38",X"E9",X"01",X"F0",X"0B",X"D5",X"C7",X"90",X"07",X"A9",X"51",X"8D",X"6C",
		X"02",X"A9",X"00",X"85",X"D4",X"20",X"0E",X"CE",X"20",X"F8",X"DE",X"50",X"08",X"A9",X"80",X"20",
		X"97",X"DD",X"4C",X"5E",X"E1",X"20",X"75",X"E2",X"A9",X"80",X"20",X"A6",X"DD",X"F0",X"03",X"4C",
		X"5E",X"E1",X"4C",X"94",X"C1",X"20",X"9C",X"E2",X"A5",X"D7",X"20",X"C8",X"D4",X"A6",X"82",X"B5",
		X"C7",X"38",X"E5",X"D4",X"B0",X"03",X"4C",X"02",X"E2",X"18",X"65",X"D7",X"90",X"03",X"69",X"01",
		X"38",X"20",X"09",X"E0",X"4C",X"38",X"E1",X"A9",X"51",X"20",X"C8",X"C1",X"A5",X"94",X"85",X"89",
		X"A5",X"95",X"85",X"8A",X"20",X"D0",X"E2",X"D0",X"01",X"60",X"20",X"F1",X"DD",X"20",X"0C",X"DE",
		X"A5",X"80",X"F0",X"0E",X"20",X"D3",X"E2",X"D0",X"06",X"20",X"1E",X"CF",X"4C",X"DA",X"D2",X"20",
		X"DA",X"D2",X"A0",X"00",X"B1",X"89",X"85",X"80",X"C8",X"B1",X"89",X"85",X"81",X"4C",X"AF",X"D0",
		X"20",X"3E",X"DE",X"A0",X"00",X"B1",X"89",X"C5",X"80",X"F0",X"01",X"60",X"C8",X"B1",X"89",X"C5",
		X"81",X"60",X"20",X"2B",X"DE",X"A0",X"02",X"A9",X"00",X"91",X"94",X"C8",X"D0",X"FB",X"20",X"04",
		X"E3",X"95",X"C1",X"A8",X"A9",X"FF",X"91",X"94",X"20",X"04",X"E3",X"90",X"F4",X"D0",X"04",X"A9",
		X"00",X"95",X"C1",X"60",X"A6",X"82",X"B5",X"C1",X"38",X"F0",X"0D",X"18",X"75",X"C7",X"90",X"0B",
		X"D0",X"06",X"A9",X"02",X"2C",X"CC",X"FE",X"60",X"69",X"01",X"38",X"60",X"20",X"D3",X"D1",X"20",
		X"CB",X"E1",X"20",X"9C",X"E2",X"20",X"7B",X"CF",X"A5",X"D6",X"85",X"87",X"A5",X"D5",X"85",X"86",
		X"A9",X"00",X"85",X"88",X"A9",X"00",X"85",X"D4",X"20",X"0E",X"CE",X"20",X"4D",X"EF",X"A4",X"82",
		X"B6",X"C7",X"CA",X"8A",X"18",X"65",X"D7",X"90",X"0C",X"E6",X"D6",X"E6",X"D6",X"D0",X"06",X"E6",
		X"D5",X"A9",X"10",X"85",X"D6",X"A5",X"87",X"18",X"69",X"02",X"20",X"E9",X"DE",X"A5",X"D5",X"C9",
		X"06",X"90",X"05",X"A9",X"52",X"20",X"C8",X"C1",X"A5",X"D6",X"38",X"E5",X"87",X"B0",X"03",X"E9",
		X"0F",X"18",X"85",X"72",X"A5",X"D5",X"E5",X"86",X"85",X"73",X"A2",X"00",X"86",X"70",X"86",X"71",
		X"AA",X"20",X"51",X"DF",X"A5",X"71",X"D0",X"07",X"A6",X"70",X"CA",X"D0",X"02",X"E6",X"88",X"CD",
		X"73",X"02",X"90",X"09",X"D0",X"CD",X"AD",X"72",X"02",X"C5",X"70",X"90",X"C6",X"A9",X"01",X"20",
		X"F6",X"D4",X"18",X"69",X"01",X"A6",X"82",X"95",X"C1",X"20",X"1E",X"F1",X"20",X"FD",X"DD",X"A5",
		X"88",X"D0",X"15",X"20",X"5E",X"DE",X"20",X"1E",X"CF",X"20",X"D0",X"D6",X"20",X"1E",X"F1",X"20",
		X"FD",X"DD",X"20",X"E2",X"E2",X"4C",X"D4",X"E3",X"20",X"1E",X"CF",X"20",X"D0",X"D6",X"20",X"E2",
		X"E2",X"20",X"19",X"DE",X"20",X"5E",X"DE",X"20",X"0C",X"DE",X"A5",X"80",X"48",X"A5",X"81",X"48",
		X"20",X"3E",X"DE",X"A5",X"81",X"48",X"A5",X"80",X"48",X"20",X"45",X"DF",X"AA",X"D0",X"0A",X"20",
		X"4E",X"E4",X"A9",X"10",X"20",X"E9",X"DE",X"E6",X"86",X"68",X"20",X"8D",X"DD",X"68",X"20",X"8D",
		X"DD",X"68",X"85",X"81",X"68",X"85",X"80",X"F0",X"0F",X"A5",X"86",X"C5",X"D5",X"D0",X"A7",X"20",
		X"45",X"DF",X"C5",X"D6",X"90",X"A0",X"F0",X"B0",X"20",X"45",X"DF",X"48",X"A9",X"00",X"20",X"DC",
		X"DE",X"A9",X"00",X"A8",X"91",X"94",X"C8",X"68",X"38",X"E9",X"01",X"91",X"94",X"20",X"6C",X"DE",
		X"20",X"99",X"D5",X"20",X"F4",X"EE",X"20",X"0E",X"CE",X"20",X"1E",X"CF",X"20",X"F8",X"DE",X"70",
		X"03",X"4C",X"75",X"E2",X"A9",X"80",X"20",X"97",X"DD",X"A9",X"50",X"20",X"C8",X"C1",X"20",X"1E",
		X"F1",X"20",X"1E",X"CF",X"20",X"F1",X"DD",X"20",X"93",X"DF",X"48",X"20",X"C1",X"DE",X"A6",X"82",
		X"B5",X"CD",X"A8",X"68",X"AA",X"A9",X"10",X"20",X"A5",X"DE",X"A9",X"00",X"20",X"DC",X"DE",X"A0",
		X"02",X"B1",X"94",X"48",X"A9",X"00",X"20",X"C8",X"D4",X"68",X"18",X"69",X"01",X"91",X"94",X"0A",
		X"69",X"04",X"85",X"89",X"A8",X"38",X"E9",X"02",X"85",X"8A",X"A5",X"80",X"85",X"87",X"91",X"94",
		X"C8",X"A5",X"81",X"85",X"88",X"91",X"94",X"A0",X"00",X"98",X"91",X"94",X"C8",X"A9",X"11",X"91",
		X"94",X"A9",X"10",X"20",X"C8",X"D4",X"20",X"50",X"DE",X"20",X"99",X"D5",X"A6",X"82",X"B5",X"CD",
		X"48",X"20",X"9E",X"DF",X"A6",X"82",X"95",X"CD",X"68",X"AE",X"57",X"02",X"95",X"A7",X"A9",X"00",
		X"20",X"C8",X"D4",X"A0",X"00",X"A5",X"80",X"91",X"94",X"C8",X"A5",X"81",X"91",X"94",X"4C",X"DE",
		X"E4",X"20",X"93",X"DF",X"A6",X"82",X"20",X"1B",X"DF",X"A9",X"00",X"20",X"C8",X"D4",X"C6",X"8A",
		X"C6",X"8A",X"A4",X"89",X"A5",X"87",X"91",X"94",X"C8",X"A5",X"88",X"91",X"94",X"20",X"5E",X"DE",
		X"20",X"99",X"D5",X"A4",X"8A",X"C0",X"03",X"B0",X"D8",X"4C",X"1E",X"CF",X"00",X"A0",X"4F",X"CB",
		X"20",X"21",X"22",X"23",X"24",X"27",X"D2",X"45",X"41",X"44",X"89",X"52",X"83",X"20",X"54",X"4F",
		X"4F",X"20",X"4C",X"41",X"52",X"47",X"C5",X"50",X"8B",X"06",X"20",X"50",X"52",X"45",X"53",X"45",
		X"4E",X"D4",X"51",X"CF",X"56",X"45",X"52",X"46",X"4C",X"4F",X"57",X"20",X"49",X"4E",X"8B",X"25",
		X"28",X"8A",X"89",X"26",X"8A",X"20",X"50",X"52",X"4F",X"54",X"45",X"43",X"54",X"20",X"4F",X"CE",
		X"29",X"88",X"20",X"49",X"44",X"85",X"30",X"31",X"32",X"33",X"34",X"D3",X"59",X"4E",X"54",X"41",
		X"58",X"89",X"60",X"8A",X"03",X"84",X"63",X"83",X"20",X"45",X"58",X"49",X"53",X"54",X"D3",X"64",
		X"83",X"20",X"54",X"59",X"50",X"45",X"85",X"65",X"CE",X"4F",X"20",X"42",X"4C",X"4F",X"43",X"CB",
		X"66",X"67",X"C9",X"4C",X"4C",X"45",X"47",X"41",X"4C",X"20",X"54",X"52",X"41",X"43",X"4B",X"20",
		X"4F",X"52",X"20",X"53",X"45",X"43",X"54",X"4F",X"D2",X"61",X"83",X"06",X"84",X"39",X"62",X"83",
		X"06",X"87",X"01",X"83",X"53",X"20",X"53",X"43",X"52",X"41",X"54",X"43",X"48",X"45",X"C4",X"70",
		X"CE",X"4F",X"20",X"43",X"48",X"41",X"4E",X"4E",X"45",X"CC",X"71",X"C4",X"49",X"52",X"89",X"72",
		X"88",X"20",X"46",X"55",X"4C",X"CC",X"73",X"CA",X"49",X"46",X"46",X"59",X"44",X"4F",X"53",X"20",
		X"35",X"2E",X"30",X"20",X"31",X"35",X"34",X"B1",X"74",X"C4",X"52",X"49",X"56",X"45",X"06",X"20",
		X"52",X"45",X"41",X"44",X"D9",X"09",X"C5",X"52",X"52",X"4F",X"D2",X"0A",X"D7",X"52",X"49",X"54",
		X"C5",X"03",X"C6",X"49",X"4C",X"C5",X"04",X"CF",X"50",X"45",X"CE",X"05",X"CD",X"49",X"53",X"4D",
		X"41",X"54",X"43",X"C8",X"06",X"CE",X"4F",X"D4",X"07",X"C6",X"4F",X"55",X"4E",X"C4",X"08",X"C4",
		X"49",X"53",X"CB",X"0B",X"D2",X"45",X"43",X"4F",X"52",X"C4",X"48",X"86",X"F9",X"8A",X"0A",X"AA",
		X"B5",X"06",X"85",X"80",X"B5",X"07",X"85",X"81",X"68",X"29",X"0F",X"F0",X"08",X"C9",X"0F",X"D0",
		X"06",X"A9",X"74",X"D0",X"08",X"A9",X"06",X"09",X"20",X"AA",X"CA",X"CA",X"8A",X"48",X"AD",X"2A",
		X"02",X"C9",X"00",X"D0",X"0F",X"A9",X"FF",X"8D",X"2A",X"02",X"68",X"20",X"C7",X"E6",X"20",X"42",
		X"D0",X"4C",X"48",X"E6",X"68",X"20",X"C7",X"E6",X"20",X"BD",X"C1",X"A9",X"00",X"8D",X"F9",X"02",
		X"20",X"2C",X"C1",X"20",X"DA",X"D4",X"A9",X"00",X"85",X"A3",X"A2",X"45",X"9A",X"A5",X"84",X"29",
		X"0F",X"85",X"83",X"C9",X"0F",X"F0",X"31",X"78",X"A5",X"79",X"D0",X"1C",X"A5",X"7A",X"D0",X"10",
		X"A6",X"83",X"BD",X"2B",X"02",X"C9",X"FF",X"F0",X"1F",X"29",X"0F",X"85",X"82",X"4C",X"8E",X"E6",
		X"20",X"EB",X"D0",X"EA",X"EA",X"EA",X"D0",X"06",X"20",X"07",X"D1",X"EA",X"EA",X"EA",X"20",X"25",
		X"D1",X"C9",X"04",X"B0",X"03",X"20",X"27",X"D2",X"4C",X"E7",X"EB",X"AA",X"A9",X"00",X"F8",X"E0",
		X"00",X"F0",X"07",X"18",X"69",X"01",X"CA",X"4C",X"9F",X"E6",X"D8",X"AA",X"4A",X"4A",X"4A",X"4A",
		X"20",X"B4",X"E6",X"8A",X"29",X"0F",X"09",X"30",X"91",X"A5",X"C8",X"60",X"20",X"23",X"C1",X"A9",
		X"00",X"A0",X"00",X"84",X"80",X"84",X"81",X"A0",X"00",X"A2",X"D5",X"86",X"A5",X"A2",X"02",X"86",
		X"A6",X"20",X"AB",X"E6",X"A9",X"2C",X"91",X"A5",X"C8",X"AD",X"D5",X"02",X"8D",X"43",X"02",X"8A",
		X"20",X"06",X"E7",X"A9",X"2C",X"91",X"A5",X"C8",X"A5",X"80",X"20",X"9B",X"E6",X"A9",X"2C",X"91",
		X"A5",X"C8",X"A5",X"81",X"20",X"9B",X"E6",X"88",X"98",X"18",X"69",X"D5",X"8D",X"49",X"02",X"E6",
		X"A5",X"A9",X"88",X"85",X"F7",X"60",X"AA",X"A5",X"86",X"48",X"A5",X"87",X"48",X"A9",X"FC",X"85",
		X"86",X"A9",X"E4",X"85",X"87",X"8A",X"A2",X"00",X"C1",X"86",X"F0",X"21",X"48",X"20",X"75",X"E7",
		X"90",X"05",X"20",X"75",X"E7",X"90",X"FB",X"A5",X"87",X"C9",X"E6",X"90",X"08",X"D0",X"0A",X"A9",
		X"0A",X"C5",X"86",X"90",X"04",X"68",X"4C",X"18",X"E7",X"68",X"4C",X"4D",X"E7",X"20",X"67",X"E7",
		X"90",X"FB",X"20",X"54",X"E7",X"20",X"67",X"E7",X"90",X"F8",X"20",X"54",X"E7",X"68",X"85",X"87",
		X"68",X"85",X"86",X"60",X"C9",X"20",X"B0",X"0B",X"AA",X"A9",X"20",X"91",X"A5",X"C8",X"8A",X"20",
		X"06",X"E7",X"60",X"91",X"A5",X"C8",X"60",X"E6",X"86",X"D0",X"02",X"E6",X"87",X"A1",X"86",X"0A",
		X"A1",X"86",X"29",X"7F",X"60",X"20",X"6D",X"E7",X"E6",X"86",X"D0",X"02",X"E6",X"87",X"60",X"60",
		X"60",X"20",X"F6",X"FE",X"0A",X"10",X"03",X"4C",X"2D",X"FF",X"20",X"25",X"D1",X"AA",X"F0",X"0C",
		X"C9",X"03",X"B0",X"08",X"AD",X"54",X"02",X"D0",X"03",X"4C",X"33",X"FB",X"38",X"66",X"98",X"4C",
		X"3B",X"FB",X"60",X"A9",X"8D",X"20",X"68",X"C2",X"20",X"58",X"F2",X"AD",X"78",X"02",X"48",X"A9",
		X"01",X"8D",X"78",X"02",X"A9",X"FF",X"85",X"86",X"20",X"4F",X"C4",X"AD",X"80",X"02",X"D0",X"05",
		X"A9",X"39",X"20",X"C8",X"C1",X"68",X"8D",X"78",X"02",X"AD",X"80",X"02",X"85",X"80",X"AD",X"85",
		X"02",X"85",X"81",X"A9",X"03",X"20",X"77",X"D4",X"A9",X"00",X"85",X"87",X"20",X"39",X"E8",X"85",
		X"88",X"20",X"4B",X"E8",X"20",X"39",X"E8",X"85",X"89",X"20",X"4B",X"E8",X"A5",X"86",X"F0",X"0A",
		X"A5",X"88",X"48",X"A5",X"89",X"48",X"A9",X"00",X"85",X"86",X"20",X"39",X"E8",X"85",X"8A",X"20",
		X"4B",X"E8",X"20",X"39",X"E8",X"A0",X"00",X"91",X"88",X"20",X"4B",X"E8",X"A5",X"88",X"18",X"69",
		X"01",X"85",X"88",X"90",X"02",X"E6",X"89",X"C6",X"8A",X"D0",X"E7",X"20",X"35",X"CA",X"A5",X"85",
		X"C5",X"87",X"F0",X"08",X"20",X"3E",X"DE",X"A9",X"50",X"20",X"45",X"E6",X"A5",X"F8",X"D0",X"A8",
		X"68",X"85",X"89",X"68",X"85",X"88",X"6C",X"88",X"00",X"20",X"35",X"CA",X"A5",X"F8",X"D0",X"08",
		X"20",X"3E",X"DE",X"A9",X"51",X"20",X"45",X"E6",X"A5",X"85",X"60",X"18",X"65",X"87",X"69",X"00",
		X"85",X"87",X"60",X"AD",X"01",X"18",X"A9",X"01",X"85",X"7C",X"60",X"78",X"A9",X"00",X"85",X"98",
		X"85",X"79",X"85",X"7A",X"85",X"7C",X"A2",X"45",X"9A",X"2C",X"00",X"18",X"10",X"5C",X"A0",X"80",
		X"84",X"F8",X"84",X"7D",X"A9",X"12",X"8D",X"00",X"18",X"20",X"F6",X"FE",X"20",X"C9",X"E9",X"D0",
		X"02",X"85",X"98",X"C9",X"3F",X"F0",X"0A",X"C9",X"5F",X"F0",X"10",X"C5",X"78",X"D0",X"06",X"84",
		X"7A",X"86",X"79",X"F0",X"30",X"C5",X"77",X"D0",X"06",X"84",X"79",X"86",X"7A",X"F0",X"26",X"C9",
		X"61",X"D0",X"08",X"A6",X"7A",X"F0",X"04",X"A9",X"60",X"85",X"98",X"AA",X"29",X"60",X"C9",X"60",
		X"D0",X"3A",X"86",X"84",X"8A",X"29",X"0F",X"85",X"83",X"8A",X"29",X"F0",X"C9",X"E0",X"D0",X"37",
		X"58",X"20",X"C0",X"DA",X"78",X"AD",X"00",X"18",X"30",X"B2",X"A2",X"00",X"86",X"7D",X"29",X"EF",
		X"8D",X"00",X"18",X"A5",X"79",X"F0",X"06",X"20",X"2E",X"EA",X"4C",X"E7",X"EB",X"A5",X"7A",X"F0",
		X"08",X"A9",X"08",X"8D",X"00",X"18",X"20",X"09",X"E9",X"4C",X"4E",X"EA",X"A5",X"79",X"05",X"7A",
		X"D0",X"05",X"A9",X"10",X"8D",X"00",X"18",X"AD",X"00",X"18",X"10",X"CE",X"30",X"F9",X"20",X"10",
		X"F9",X"4C",X"18",X"F4",X"0A",X"0A",X"0B",X"0C",X"F9",X"78",X"20",X"EB",X"D0",X"B0",X"5D",X"A5",
		X"98",X"F0",X"05",X"A2",X"46",X"4C",X"81",X"E7",X"A6",X"82",X"B4",X"F2",X"10",X"4E",X"AD",X"00",
		X"18",X"29",X"F7",X"8D",X"00",X"18",X"4A",X"90",X"08",X"20",X"6D",X"E9",X"98",X"29",X"08",X"D0",
		X"03",X"20",X"66",X"E9",X"20",X"AE",X"E9",X"20",X"6D",X"E9",X"A0",X"08",X"A6",X"82",X"7E",X"3E",
		X"02",X"20",X"9C",X"E9",X"B0",X"02",X"09",X"02",X"20",X"A1",X"E9",X"20",X"BA",X"E9",X"A2",X"0B",
		X"CA",X"D0",X"FD",X"09",X"08",X"20",X"9F",X"E9",X"88",X"D0",X"E1",X"20",X"66",X"E9",X"58",X"20",
		X"AA",X"D3",X"78",X"4C",X"18",X"E9",X"20",X"59",X"EA",X"6A",X"90",X"FA",X"60",X"20",X"59",X"EA",
		X"6A",X"B0",X"FA",X"60",X"A1",X"99",X"85",X"80",X"F6",X"99",X"A1",X"99",X"85",X"81",X"20",X"64",
		X"FB",X"20",X"D3",X"D0",X"20",X"A4",X"D0",X"A6",X"80",X"D0",X"03",X"99",X"44",X"02",X"60",X"F0",
		X"F6",X"58",X"20",X"AA",X"D3",X"78",X"4C",X"0F",X"E9",X"4C",X"4E",X"EA",X"AD",X"00",X"18",X"29",
		X"FD",X"8D",X"00",X"18",X"60",X"AD",X"00",X"18",X"09",X"02",X"8D",X"00",X"18",X"60",X"AD",X"00",
		X"18",X"09",X"08",X"8D",X"00",X"18",X"60",X"AD",X"00",X"18",X"29",X"F7",X"8D",X"00",X"18",X"60",
		X"AD",X"00",X"18",X"CD",X"00",X"18",X"D0",X"F8",X"60",X"A9",X"08",X"85",X"4B",X"20",X"17",X"EA",
		X"D0",X"FB",X"20",X"9C",X"E9",X"20",X"20",X"FF",X"A2",X"90",X"20",X"17",X"EA",X"D0",X"0D",X"CA",
		X"30",X"F8",X"20",X"83",X"F6",X"86",X"F8",X"20",X"17",X"EA",X"F0",X"FB",X"A2",X"0C",X"AD",X"00",
		X"18",X"85",X"44",X"29",X"04",X"F0",X"08",X"CA",X"D0",X"F4",X"20",X"74",X"F6",X"F0",X"EF",X"A5",
		X"44",X"49",X"01",X"4A",X"66",X"85",X"20",X"17",X"EA",X"F0",X"FB",X"C6",X"4B",X"D0",X"DD",X"20",
		X"A5",X"E9",X"A2",X"00",X"A5",X"85",X"60",X"20",X"59",X"EA",X"29",X"04",X"60",X"0F",X"07",X"0D",
		X"05",X"0B",X"03",X"09",X"01",X"0E",X"06",X"0C",X"04",X"0A",X"02",X"08",X"00",X"60",X"78",X"20",
		X"07",X"D1",X"B0",X"05",X"B5",X"F2",X"6A",X"B0",X"0B",X"A5",X"84",X"29",X"F0",X"C9",X"F0",X"F0",
		X"03",X"4C",X"4E",X"EA",X"20",X"C1",X"FB",X"EA",X"20",X"69",X"F7",X"4C",X"2E",X"EA",X"A9",X"00",
		X"8D",X"00",X"18",X"4C",X"E7",X"EB",X"4C",X"5B",X"E8",X"A5",X"7D",X"F0",X"06",X"AD",X"00",X"18",
		X"10",X"09",X"60",X"AD",X"00",X"18",X"10",X"FA",X"4C",X"5B",X"E8",X"4C",X"CA",X"E8",X"A2",X"00",
		X"2C",X"A6",X"6F",X"9A",X"BA",X"A9",X"08",X"0D",X"00",X"1C",X"4C",X"EA",X"FE",X"98",X"18",X"69",
		X"01",X"D0",X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"1C",X"29",X"F7",X"8D",X"00",X"1C",X"98",X"18",
		X"69",X"01",X"D0",X"FC",X"88",X"D0",X"F8",X"CA",X"10",X"DB",X"E0",X"FC",X"D0",X"F0",X"F0",X"D4",
		X"78",X"D8",X"A2",X"FF",X"4C",X"10",X"FF",X"E8",X"A0",X"00",X"A2",X"00",X"8A",X"95",X"00",X"E8",
		X"D0",X"FA",X"8A",X"D5",X"00",X"D0",X"B7",X"F6",X"00",X"C8",X"D0",X"FB",X"D5",X"00",X"D0",X"AE",
		X"94",X"00",X"B5",X"00",X"D0",X"A8",X"E8",X"D0",X"E9",X"E6",X"6F",X"86",X"76",X"A9",X"00",X"85",
		X"75",X"A8",X"A2",X"20",X"18",X"C6",X"76",X"71",X"75",X"C8",X"D0",X"FB",X"CA",X"D0",X"F6",X"69",
		X"00",X"AA",X"C5",X"76",X"D0",X"39",X"E0",X"C0",X"D0",X"DF",X"A9",X"01",X"85",X"76",X"E6",X"6F",
		X"A2",X"07",X"98",X"18",X"65",X"76",X"91",X"75",X"C8",X"D0",X"F7",X"E6",X"76",X"CA",X"D0",X"F2",
		X"A2",X"07",X"C6",X"76",X"88",X"98",X"18",X"65",X"76",X"D1",X"75",X"D0",X"12",X"49",X"FF",X"91",
		X"75",X"51",X"75",X"91",X"75",X"D0",X"08",X"98",X"D0",X"EA",X"CA",X"D0",X"E5",X"F0",X"03",X"4C",
		X"71",X"EA",X"A2",X"45",X"9A",X"AD",X"00",X"1C",X"29",X"F7",X"8D",X"00",X"1C",X"A9",X"01",X"8D",
		X"0C",X"18",X"A9",X"82",X"8D",X"0D",X"18",X"8D",X"0E",X"18",X"AD",X"00",X"18",X"29",X"60",X"0A",
		X"2A",X"2A",X"2A",X"09",X"48",X"85",X"78",X"49",X"60",X"85",X"77",X"A2",X"00",X"A0",X"00",X"A9",
		X"00",X"95",X"99",X"E8",X"B9",X"E0",X"FE",X"95",X"99",X"E8",X"C8",X"C0",X"05",X"D0",X"F0",X"A9",
		X"00",X"95",X"99",X"E8",X"A9",X"02",X"95",X"99",X"E8",X"A9",X"D5",X"95",X"99",X"E8",X"A9",X"02",
		X"95",X"99",X"A9",X"FF",X"A2",X"12",X"9D",X"2B",X"02",X"CA",X"10",X"FA",X"A2",X"05",X"95",X"A7",
		X"95",X"AE",X"95",X"CD",X"CA",X"10",X"F7",X"A9",X"05",X"85",X"AB",X"A9",X"06",X"85",X"AC",X"A9",
		X"FF",X"85",X"AD",X"85",X"B4",X"A9",X"05",X"8D",X"3B",X"02",X"A9",X"84",X"8D",X"3A",X"02",X"A9",
		X"0F",X"8D",X"56",X"02",X"A9",X"01",X"85",X"F6",X"A9",X"88",X"85",X"F7",X"A9",X"E0",X"8D",X"4F",
		X"02",X"A9",X"FF",X"8D",X"50",X"02",X"A9",X"01",X"85",X"1C",X"85",X"1D",X"20",X"63",X"CB",X"20",
		X"FA",X"CE",X"20",X"59",X"F2",X"A9",X"22",X"85",X"65",X"A9",X"EB",X"85",X"66",X"A9",X"00",X"85",
		X"69",X"A9",X"05",X"85",X"6A",X"A9",X"73",X"20",X"C1",X"E6",X"A9",X"00",X"8D",X"00",X"18",X"A9",
		X"1A",X"8D",X"02",X"18",X"20",X"80",X"E7",X"58",X"AD",X"00",X"18",X"29",X"E5",X"8D",X"00",X"18",
		X"AD",X"55",X"02",X"F0",X"0A",X"A9",X"00",X"8D",X"55",X"02",X"85",X"67",X"20",X"46",X"C1",X"58",
		X"A5",X"7C",X"F0",X"03",X"4C",X"5B",X"E8",X"58",X"A9",X"0E",X"85",X"72",X"A9",X"00",X"85",X"6F",
		X"85",X"70",X"A6",X"72",X"BD",X"2B",X"02",X"C9",X"FF",X"F0",X"10",X"29",X"3F",X"85",X"82",X"20",
		X"93",X"DF",X"AA",X"BD",X"5B",X"02",X"29",X"01",X"AA",X"F6",X"6F",X"C6",X"72",X"10",X"E3",X"A0",
		X"04",X"B9",X"00",X"00",X"10",X"05",X"29",X"01",X"AA",X"F6",X"6F",X"88",X"10",X"F3",X"78",X"AD",
		X"00",X"1C",X"29",X"F7",X"48",X"A5",X"7F",X"85",X"86",X"A9",X"00",X"85",X"7F",X"A5",X"6F",X"F0",
		X"0B",X"A5",X"1C",X"F0",X"03",X"20",X"13",X"D3",X"68",X"09",X"08",X"48",X"E6",X"7F",X"A5",X"70",
		X"F0",X"0B",X"A5",X"1D",X"F0",X"03",X"20",X"13",X"D3",X"68",X"09",X"00",X"48",X"A5",X"86",X"85",
		X"7F",X"68",X"AE",X"6C",X"02",X"F0",X"21",X"AD",X"00",X"1C",X"E0",X"80",X"D0",X"03",X"4C",X"8B",
		X"EC",X"AE",X"05",X"18",X"30",X"12",X"A2",X"A0",X"8E",X"05",X"18",X"CE",X"6C",X"02",X"D0",X"08",
		X"4D",X"6D",X"02",X"A2",X"10",X"8E",X"6C",X"02",X"8D",X"00",X"1C",X"4C",X"FF",X"EB",X"A9",X"00",
		X"85",X"83",X"A9",X"01",X"20",X"E2",X"D1",X"A9",X"00",X"20",X"C8",X"D4",X"A6",X"82",X"A9",X"00",
		X"9D",X"44",X"02",X"20",X"93",X"DF",X"AA",X"A5",X"7F",X"9D",X"5B",X"02",X"A9",X"01",X"20",X"F1",
		X"CF",X"A9",X"04",X"20",X"F1",X"CF",X"A9",X"01",X"20",X"F1",X"CF",X"20",X"F1",X"CF",X"AD",X"72",
		X"02",X"20",X"F1",X"CF",X"A9",X"00",X"20",X"F1",X"CF",X"20",X"59",X"ED",X"20",X"93",X"DF",X"0A",
		X"AA",X"D6",X"99",X"D6",X"99",X"A9",X"00",X"20",X"F1",X"CF",X"A9",X"01",X"20",X"F1",X"CF",X"20",
		X"F1",X"CF",X"20",X"CE",X"C6",X"90",X"2C",X"AD",X"72",X"02",X"20",X"F1",X"CF",X"AD",X"73",X"02",
		X"20",X"F1",X"CF",X"20",X"59",X"ED",X"A9",X"00",X"20",X"F1",X"CF",X"D0",X"DD",X"20",X"93",X"DF",
		X"0A",X"AA",X"A9",X"00",X"95",X"99",X"A9",X"88",X"A4",X"82",X"8D",X"54",X"02",X"99",X"F2",X"00",
		X"A5",X"85",X"60",X"AD",X"72",X"02",X"20",X"F1",X"CF",X"AD",X"73",X"02",X"20",X"F1",X"CF",X"20",
		X"59",X"ED",X"20",X"93",X"DF",X"0A",X"AA",X"D6",X"99",X"D6",X"99",X"A9",X"00",X"20",X"F1",X"CF",
		X"20",X"F1",X"CF",X"20",X"F1",X"CF",X"20",X"93",X"DF",X"0A",X"A8",X"B9",X"99",X"00",X"A6",X"82",
		X"9D",X"44",X"02",X"DE",X"44",X"02",X"4C",X"0D",X"ED",X"A0",X"00",X"B9",X"B1",X"02",X"20",X"F1",
		X"CF",X"C8",X"C0",X"1B",X"D0",X"F5",X"60",X"20",X"37",X"D1",X"F0",X"01",X"60",X"85",X"85",X"A4",
		X"82",X"B9",X"44",X"02",X"F0",X"08",X"A9",X"80",X"99",X"F2",X"00",X"A5",X"85",X"60",X"48",X"20",
		X"EA",X"EC",X"68",X"60",X"20",X"D1",X"C1",X"20",X"42",X"D0",X"A9",X"40",X"8D",X"F9",X"02",X"20",
		X"B7",X"EE",X"A9",X"00",X"8D",X"92",X"02",X"20",X"AC",X"C5",X"D0",X"3D",X"A9",X"00",X"85",X"81",
		X"AD",X"85",X"FE",X"85",X"80",X"20",X"E5",X"ED",X"A9",X"00",X"8D",X"F9",X"02",X"20",X"FF",X"EE",
		X"4C",X"94",X"C1",X"C8",X"B1",X"94",X"48",X"C8",X"B1",X"94",X"48",X"A0",X"13",X"B1",X"94",X"F0",
		X"0A",X"85",X"80",X"C8",X"B1",X"94",X"85",X"81",X"20",X"E5",X"ED",X"68",X"85",X"81",X"68",X"85",
		X"80",X"20",X"E5",X"ED",X"20",X"04",X"C6",X"F0",X"C3",X"A0",X"00",X"B1",X"94",X"30",X"D4",X"20",
		X"B6",X"C8",X"4C",X"D4",X"ED",X"20",X"5F",X"D5",X"20",X"90",X"EF",X"20",X"75",X"D4",X"A9",X"00",
		X"20",X"C8",X"D4",X"20",X"A4",X"D0",X"A5",X"80",X"D0",X"03",X"4C",X"27",X"D2",X"20",X"90",X"EF",
		X"78",X"20",X"64",X"FB",X"58",X"4C",X"EE",X"ED",X"4D",X"D4",X"4C",X"EE",X"ED",X"20",X"12",X"C3",
		X"A5",X"E2",X"10",X"05",X"A9",X"33",X"4C",X"C8",X"C1",X"29",X"01",X"85",X"7F",X"20",X"00",X"C1",
		X"A5",X"7F",X"0A",X"AA",X"AC",X"7B",X"02",X"CC",X"74",X"02",X"F0",X"1A",X"B9",X"00",X"02",X"95",
		X"12",X"B9",X"01",X"02",X"95",X"13",X"20",X"07",X"D3",X"A9",X"01",X"85",X"80",X"20",X"C6",X"C8",
		X"20",X"05",X"F0",X"4C",X"56",X"EE",X"20",X"42",X"D0",X"A6",X"7F",X"BD",X"01",X"01",X"CD",X"D5",
		X"FE",X"F0",X"03",X"4C",X"72",X"D5",X"20",X"B7",X"EE",X"A5",X"F9",X"A8",X"0A",X"AA",X"AD",X"88",
		X"FE",X"95",X"99",X"AE",X"7A",X"02",X"A9",X"1B",X"20",X"6E",X"C6",X"A0",X"12",X"A6",X"7F",X"AD",
		X"D5",X"FE",X"9D",X"01",X"01",X"8A",X"0A",X"AA",X"B5",X"12",X"91",X"94",X"C8",X"B5",X"13",X"91",
		X"94",X"C8",X"C8",X"A9",X"32",X"91",X"94",X"C8",X"AD",X"D5",X"FE",X"91",X"94",X"A0",X"02",X"91",
		X"6D",X"AD",X"85",X"FE",X"85",X"80",X"20",X"93",X"EF",X"A9",X"01",X"85",X"81",X"20",X"93",X"EF",
		X"20",X"FF",X"EE",X"20",X"05",X"F0",X"A0",X"01",X"A9",X"FF",X"91",X"6D",X"20",X"64",X"D4",X"C6",
		X"81",X"20",X"60",X"D4",X"4C",X"94",X"C1",X"20",X"D1",X"F0",X"A0",X"00",X"A9",X"12",X"91",X"6D",
		X"C8",X"98",X"91",X"6D",X"C8",X"C8",X"C8",X"A9",X"00",X"85",X"6F",X"85",X"70",X"85",X"71",X"98",
		X"4A",X"4A",X"20",X"4B",X"F2",X"91",X"6D",X"C8",X"AA",X"38",X"26",X"6F",X"26",X"70",X"26",X"71",
		X"CA",X"D0",X"F6",X"B5",X"6F",X"91",X"6D",X"C8",X"E8",X"E0",X"03",X"90",X"F6",X"C0",X"90",X"90",
		X"D6",X"4C",X"75",X"D0",X"20",X"93",X"DF",X"AA",X"BD",X"5B",X"02",X"29",X"01",X"85",X"7F",X"A4",
		X"7F",X"B9",X"51",X"02",X"D0",X"01",X"60",X"A9",X"00",X"99",X"51",X"02",X"20",X"3A",X"EF",X"A5",
		X"7F",X"0A",X"48",X"20",X"A5",X"F0",X"68",X"18",X"69",X"01",X"20",X"A5",X"F0",X"A5",X"80",X"48",
		X"A9",X"01",X"85",X"80",X"0A",X"0A",X"85",X"6D",X"20",X"20",X"F2",X"E6",X"80",X"A5",X"80",X"CD",
		X"D7",X"FE",X"90",X"F0",X"68",X"85",X"80",X"4C",X"8A",X"D5",X"20",X"0F",X"F1",X"AA",X"20",X"DF",
		X"F0",X"A6",X"F9",X"BD",X"E0",X"FE",X"85",X"6E",X"A9",X"00",X"85",X"6D",X"60",X"A6",X"7F",X"BD",
		X"FA",X"02",X"8D",X"72",X"02",X"BD",X"FC",X"02",X"8D",X"73",X"02",X"60",X"20",X"F1",X"EF",X"20",
		X"CF",X"EF",X"D0",X"21",X"B1",X"6D",X"1D",X"E9",X"EF",X"91",X"6D",X"20",X"88",X"EF",X"A4",X"6F",
		X"18",X"B1",X"6D",X"69",X"01",X"91",X"6D",X"A5",X"80",X"C9",X"12",X"F0",X"3D",X"FE",X"FA",X"02",
		X"D0",X"03",X"FE",X"FC",X"02",X"4C",X"D9",X"F7",X"A6",X"7F",X"A9",X"01",X"9D",X"51",X"02",X"60",
		X"20",X"F1",X"EF",X"20",X"CF",X"EF",X"F0",X"36",X"B1",X"6D",X"5D",X"E9",X"EF",X"91",X"6D",X"20",
		X"88",X"EF",X"A4",X"6F",X"B1",X"6D",X"38",X"E9",X"01",X"91",X"6D",X"A5",X"80",X"CD",X"85",X"FE",
		X"F0",X"0B",X"BD",X"FA",X"02",X"D0",X"03",X"DE",X"FC",X"02",X"DE",X"FA",X"02",X"BD",X"FC",X"02",
		X"D0",X"0C",X"BD",X"FA",X"02",X"C9",X"03",X"B0",X"05",X"A9",X"72",X"20",X"C7",X"E6",X"60",X"20",
		X"11",X"F0",X"98",X"85",X"6F",X"A5",X"81",X"4A",X"4A",X"4A",X"38",X"65",X"6F",X"A8",X"A5",X"81",
		X"29",X"07",X"AA",X"B1",X"6D",X"3D",X"E9",X"EF",X"60",X"01",X"02",X"04",X"08",X"10",X"20",X"40",
		X"80",X"A9",X"FF",X"2C",X"F9",X"02",X"F0",X"0C",X"10",X"0A",X"70",X"08",X"A9",X"00",X"8D",X"F9",
		X"02",X"4C",X"8A",X"D5",X"60",X"20",X"3A",X"EF",X"A0",X"00",X"98",X"91",X"6D",X"C8",X"D0",X"FB",
		X"60",X"A5",X"6F",X"48",X"A5",X"70",X"48",X"A6",X"7F",X"B5",X"FF",X"F0",X"05",X"A9",X"74",X"20",
		X"48",X"E6",X"20",X"0F",X"F1",X"85",X"6F",X"8A",X"0A",X"85",X"70",X"AA",X"A5",X"80",X"DD",X"9D",
		X"02",X"F0",X"0B",X"E8",X"86",X"70",X"DD",X"9D",X"02",X"F0",X"03",X"20",X"5B",X"F0",X"A5",X"70",
		X"A6",X"7F",X"9D",X"9B",X"02",X"0A",X"0A",X"18",X"69",X"A1",X"85",X"6D",X"A9",X"02",X"69",X"00",
		X"85",X"6E",X"A0",X"00",X"68",X"85",X"70",X"68",X"85",X"6F",X"60",X"A6",X"6F",X"20",X"DF",X"F0",
		X"A5",X"7F",X"AA",X"0A",X"1D",X"9B",X"02",X"49",X"01",X"29",X"03",X"85",X"70",X"20",X"A5",X"F0",
		X"A5",X"F9",X"0A",X"AA",X"A5",X"80",X"0A",X"0A",X"95",X"99",X"A5",X"70",X"0A",X"0A",X"A8",X"A1",
		X"99",X"99",X"A1",X"02",X"A9",X"00",X"81",X"99",X"F6",X"99",X"C8",X"98",X"29",X"03",X"D0",X"EF",
		X"A6",X"70",X"A5",X"80",X"9D",X"9D",X"02",X"AD",X"F9",X"02",X"D0",X"03",X"4C",X"8A",X"D5",X"09",
		X"80",X"8D",X"F9",X"02",X"60",X"A8",X"B9",X"9D",X"02",X"F0",X"25",X"48",X"A9",X"00",X"99",X"9D",
		X"02",X"A5",X"F9",X"0A",X"AA",X"68",X"0A",X"0A",X"95",X"99",X"98",X"0A",X"0A",X"A8",X"B9",X"A1",
		X"02",X"81",X"99",X"A9",X"00",X"99",X"A1",X"02",X"F6",X"99",X"C8",X"98",X"29",X"03",X"D0",X"EE",
		X"60",X"A5",X"7F",X"0A",X"AA",X"A9",X"00",X"9D",X"9D",X"02",X"E8",X"9D",X"9D",X"02",X"60",X"B5",
		X"A7",X"C9",X"FF",X"D0",X"25",X"8A",X"48",X"20",X"8E",X"D2",X"AA",X"10",X"05",X"A9",X"70",X"20",
		X"C8",X"C1",X"86",X"F9",X"68",X"A8",X"8A",X"09",X"80",X"99",X"A7",X"00",X"0A",X"AA",X"AD",X"85",
		X"FE",X"95",X"06",X"A9",X"00",X"95",X"07",X"4C",X"86",X"D5",X"29",X"0F",X"85",X"F9",X"60",X"A9",
		X"06",X"A6",X"7F",X"D0",X"03",X"18",X"69",X"07",X"60",X"20",X"0F",X"F1",X"AA",X"60",X"20",X"3E",
		X"DE",X"A9",X"03",X"85",X"6F",X"A9",X"01",X"0D",X"F9",X"02",X"8D",X"F9",X"02",X"20",X"11",X"F0",
		X"B1",X"6D",X"D0",X"3F",X"A5",X"81",X"85",X"81",X"A2",X"12",X"E4",X"80",X"F0",X"1C",X"B0",X"11",
		X"E6",X"80",X"A5",X"80",X"C9",X"24",X"D0",X"E5",X"CA",X"86",X"80",X"C6",X"6F",X"D0",X"DE",X"F0",
		X"09",X"C6",X"80",X"D0",X"D8",X"E8",X"D0",X"F1",X"EA",X"EA",X"A9",X"72",X"20",X"C8",X"C1",X"20",
		X"25",X"D1",X"A8",X"A5",X"80",X"20",X"4B",X"F2",X"A9",X"06",X"EA",X"C0",X"02",X"F0",X"09",X"BD",
		X"04",X"E9",X"2C",X"A5",X"69",X"AA",X"F0",X"E7",X"18",X"65",X"81",X"85",X"81",X"A5",X"80",X"20",
		X"4B",X"F2",X"8D",X"4E",X"02",X"8D",X"4D",X"02",X"C5",X"81",X"B0",X"09",X"38",X"A5",X"81",X"ED",
		X"4E",X"02",X"85",X"81",X"EA",X"20",X"FA",X"F1",X"F0",X"03",X"4C",X"90",X"EF",X"A9",X"00",X"85",
		X"81",X"20",X"FA",X"F1",X"D0",X"F4",X"4C",X"F5",X"F1",X"A9",X"01",X"0D",X"F9",X"02",X"8D",X"F9",
		X"02",X"A5",X"86",X"48",X"A9",X"01",X"85",X"86",X"AD",X"85",X"FE",X"38",X"E5",X"86",X"85",X"80",
		X"90",X"09",X"F0",X"07",X"20",X"11",X"F0",X"B1",X"6D",X"D0",X"1B",X"AD",X"85",X"FE",X"18",X"65",
		X"86",X"85",X"80",X"E6",X"86",X"CD",X"D7",X"FE",X"90",X"05",X"A9",X"67",X"20",X"45",X"E6",X"20",
		X"11",X"F0",X"B1",X"6D",X"F0",X"D2",X"68",X"85",X"86",X"A9",X"00",X"85",X"81",X"20",X"FA",X"F1",
		X"F0",X"03",X"4C",X"90",X"EF",X"A9",X"71",X"20",X"45",X"E6",X"20",X"11",X"F0",X"98",X"48",X"20",
		X"20",X"F2",X"A5",X"80",X"20",X"4B",X"F2",X"8D",X"4E",X"02",X"68",X"85",X"6F",X"A5",X"81",X"CD",
		X"4E",X"02",X"B0",X"09",X"20",X"D5",X"EF",X"D0",X"06",X"E6",X"81",X"D0",X"F0",X"A9",X"00",X"60",
		X"A5",X"6F",X"48",X"A9",X"00",X"85",X"6F",X"AC",X"86",X"FE",X"88",X"A2",X"07",X"B1",X"6D",X"3D",
		X"E9",X"EF",X"F0",X"02",X"E6",X"6F",X"CA",X"10",X"F4",X"88",X"D0",X"EF",X"B1",X"6D",X"C5",X"6F",
		X"D0",X"04",X"68",X"85",X"6F",X"60",X"A9",X"71",X"20",X"45",X"E6",X"AE",X"D6",X"FE",X"DD",X"D6",
		X"FE",X"CA",X"B0",X"FA",X"BD",X"D1",X"FE",X"60",X"60",X"A9",X"6F",X"8D",X"02",X"1C",X"29",X"F0",
		X"8D",X"00",X"1C",X"AD",X"0C",X"1C",X"29",X"FE",X"09",X"0E",X"09",X"E0",X"8D",X"0C",X"1C",X"A9",
		X"41",X"8D",X"0B",X"1C",X"A9",X"00",X"8D",X"06",X"1C",X"A9",X"3A",X"8D",X"07",X"1C",X"8D",X"05",
		X"1C",X"A9",X"7F",X"8D",X"0E",X"1C",X"A9",X"C0",X"8D",X"0D",X"1C",X"8D",X"0E",X"1C",X"A9",X"FF",
		X"85",X"3E",X"85",X"51",X"A9",X"08",X"85",X"39",X"A9",X"07",X"85",X"47",X"A9",X"05",X"85",X"62",
		X"A9",X"FA",X"85",X"63",X"A9",X"C8",X"85",X"64",X"A9",X"04",X"85",X"5E",X"A9",X"04",X"85",X"5F",
		X"BA",X"86",X"49",X"AD",X"04",X"1C",X"AD",X"0C",X"1C",X"09",X"0E",X"8D",X"0C",X"1C",X"A0",X"05",
		X"B9",X"00",X"00",X"10",X"2E",X"C9",X"D0",X"D0",X"04",X"98",X"4C",X"70",X"F3",X"29",X"01",X"F0",
		X"07",X"84",X"3F",X"A9",X"0F",X"4C",X"69",X"F9",X"AA",X"85",X"3D",X"C5",X"3E",X"F0",X"0A",X"20",
		X"7E",X"F9",X"A5",X"3D",X"85",X"3E",X"4C",X"9C",X"F9",X"A5",X"20",X"30",X"03",X"0A",X"10",X"09",
		X"4C",X"9C",X"F9",X"88",X"10",X"CA",X"4C",X"9C",X"F9",X"A9",X"20",X"85",X"20",X"A0",X"05",X"84",
		X"3F",X"20",X"93",X"F3",X"30",X"1A",X"C6",X"3F",X"10",X"F7",X"A4",X"41",X"20",X"95",X"F3",X"A5",
		X"42",X"85",X"4A",X"06",X"4A",X"A9",X"60",X"85",X"20",X"B1",X"32",X"85",X"22",X"4C",X"9C",X"F9",
		X"29",X"01",X"C5",X"3D",X"D0",X"E0",X"A5",X"22",X"F0",X"12",X"38",X"F1",X"32",X"F0",X"0D",X"49",
		X"FF",X"85",X"42",X"E6",X"42",X"A5",X"3F",X"85",X"41",X"4C",X"81",X"F3",X"A2",X"04",X"B1",X"32",
		X"85",X"40",X"DD",X"D6",X"FE",X"CA",X"B0",X"FA",X"BD",X"D1",X"FE",X"85",X"43",X"8A",X"0A",X"0A",
		X"0A",X"0A",X"0A",X"85",X"44",X"AD",X"00",X"1C",X"29",X"9F",X"05",X"44",X"20",X"E4",X"FA",X"A6",
		X"3D",X"A5",X"45",X"C9",X"40",X"F0",X"15",X"C9",X"60",X"F0",X"03",X"4C",X"B1",X"F3",X"A5",X"3F",
		X"18",X"69",X"03",X"85",X"31",X"A9",X"00",X"85",X"30",X"6C",X"30",X"00",X"20",X"D3",X"FA",X"D0",
		X"0F",X"A9",X"13",X"8D",X"07",X"1C",X"4C",X"06",X"F3",X"A4",X"85",X"4A",X"A9",X"01",X"85",X"22",
		X"4C",X"69",X"F9",X"A4",X"3F",X"B9",X"00",X"00",X"48",X"10",X"10",X"29",X"78",X"85",X"45",X"98",
		X"0A",X"69",X"06",X"85",X"32",X"98",X"18",X"69",X"03",X"85",X"31",X"A0",X"00",X"84",X"30",X"68",
		X"60",X"A2",X"5A",X"86",X"4B",X"A2",X"00",X"A9",X"52",X"85",X"24",X"20",X"56",X"F5",X"50",X"FE",
		X"B8",X"AD",X"01",X"1C",X"C5",X"24",X"D0",X"3F",X"50",X"FE",X"B8",X"AD",X"01",X"1C",X"95",X"25",
		X"E8",X"E0",X"07",X"D0",X"F3",X"20",X"97",X"F4",X"A0",X"04",X"A9",X"00",X"59",X"16",X"00",X"88",
		X"10",X"FA",X"C9",X"00",X"D0",X"38",X"A6",X"3E",X"A5",X"18",X"95",X"22",X"A5",X"45",X"C9",X"30",
		X"F0",X"1E",X"A5",X"3E",X"0A",X"A8",X"B9",X"12",X"00",X"C5",X"16",X"D0",X"1E",X"B9",X"13",X"00",
		X"C5",X"17",X"D0",X"17",X"4C",X"23",X"F4",X"C6",X"4B",X"D0",X"B0",X"A9",X"02",X"20",X"69",X"F9",
		X"A5",X"16",X"85",X"12",X"A5",X"17",X"85",X"13",X"A9",X"01",X"2C",X"A9",X"0B",X"2C",X"A9",X"09",
		X"4C",X"69",X"F9",X"A9",X"7F",X"85",X"4C",X"A5",X"19",X"18",X"69",X"02",X"C5",X"43",X"90",X"02",
		X"E5",X"43",X"85",X"4D",X"A2",X"05",X"86",X"3F",X"A2",X"FF",X"20",X"93",X"F3",X"10",X"44",X"85",
		X"44",X"29",X"01",X"C5",X"3E",X"D0",X"3C",X"A0",X"00",X"B1",X"32",X"C5",X"40",X"D0",X"34",X"A5",
		X"45",X"C9",X"60",X"F0",X"0C",X"A0",X"01",X"38",X"B1",X"32",X"E5",X"4D",X"10",X"03",X"18",X"65",
		X"43",X"C5",X"4C",X"B0",X"1E",X"48",X"A5",X"45",X"F0",X"14",X"68",X"C9",X"09",X"90",X"14",X"C9",
		X"0C",X"B0",X"10",X"85",X"4C",X"A5",X"3F",X"AA",X"69",X"03",X"85",X"31",X"D0",X"05",X"68",X"C9",
		X"06",X"90",X"F0",X"C6",X"3F",X"10",X"B3",X"8A",X"10",X"03",X"4C",X"9C",X"F9",X"86",X"3F",X"20",
		X"93",X"F3",X"A5",X"45",X"4C",X"CA",X"F4",X"A5",X"30",X"48",X"A5",X"31",X"48",X"A9",X"24",X"85",
		X"30",X"A9",X"00",X"85",X"31",X"A9",X"00",X"85",X"34",X"20",X"E6",X"F7",X"A5",X"55",X"85",X"18",
		X"A5",X"54",X"85",X"19",X"A5",X"53",X"85",X"1A",X"20",X"E6",X"F7",X"A5",X"52",X"85",X"17",X"A5",
		X"53",X"85",X"16",X"68",X"85",X"31",X"68",X"85",X"30",X"60",X"C9",X"00",X"F0",X"03",X"4C",X"6E",
		X"F5",X"20",X"0A",X"F5",X"50",X"FE",X"B8",X"AD",X"01",X"1C",X"91",X"30",X"C8",X"D0",X"F5",X"A0",
		X"BA",X"50",X"FE",X"B8",X"AD",X"01",X"1C",X"99",X"00",X"01",X"C8",X"D0",X"F4",X"20",X"E0",X"F8",
		X"A5",X"38",X"C5",X"47",X"F0",X"05",X"A9",X"04",X"4C",X"69",X"F9",X"A5",X"4B",X"EA",X"C5",X"3A",
		X"F0",X"03",X"A9",X"05",X"2C",X"A9",X"01",X"4C",X"69",X"F9",X"20",X"10",X"F5",X"4C",X"56",X"F5",
		X"A5",X"3D",X"0A",X"AA",X"B5",X"12",X"85",X"16",X"B5",X"13",X"85",X"17",X"A0",X"00",X"B1",X"32",
		X"85",X"18",X"C8",X"B1",X"32",X"85",X"19",X"A9",X"00",X"45",X"16",X"45",X"17",X"45",X"18",X"45",
		X"19",X"85",X"1A",X"20",X"34",X"F9",X"A2",X"5A",X"20",X"56",X"F5",X"A0",X"00",X"50",X"FE",X"B8",
		X"AD",X"01",X"1C",X"D9",X"24",X"00",X"D0",X"06",X"C8",X"C0",X"08",X"D0",X"F0",X"60",X"CA",X"D0",
		X"E7",X"A9",X"02",X"4C",X"69",X"F9",X"A9",X"D0",X"8D",X"05",X"18",X"A9",X"03",X"2C",X"05",X"18",
		X"10",X"F1",X"2C",X"00",X"1C",X"30",X"F6",X"AD",X"01",X"1C",X"B8",X"A0",X"00",X"60",X"C9",X"10",
		X"F0",X"03",X"4C",X"91",X"F6",X"20",X"E9",X"F5",X"85",X"3A",X"AD",X"00",X"1C",X"29",X"10",X"D0",
		X"05",X"A9",X"08",X"4C",X"69",X"F9",X"20",X"8F",X"F7",X"20",X"10",X"F5",X"A2",X"09",X"50",X"FE",
		X"B8",X"CA",X"D0",X"FA",X"A9",X"FF",X"8D",X"03",X"1C",X"AD",X"0C",X"1C",X"29",X"1F",X"09",X"C0",
		X"8D",X"0C",X"1C",X"A9",X"FF",X"A2",X"05",X"8D",X"01",X"1C",X"B8",X"50",X"FE",X"B8",X"CA",X"D0",
		X"FA",X"A0",X"BB",X"B9",X"00",X"01",X"50",X"FE",X"B8",X"8D",X"01",X"1C",X"C8",X"D0",X"F4",X"B1",
		X"30",X"50",X"FE",X"B8",X"8D",X"01",X"1C",X"C8",X"D0",X"F5",X"50",X"FE",X"AD",X"0C",X"1C",X"09",
		X"E0",X"8D",X"0C",X"1C",X"A9",X"00",X"8D",X"03",X"1C",X"20",X"0D",X"F9",X"A4",X"3F",X"B9",X"00",
		X"00",X"49",X"30",X"99",X"00",X"00",X"4C",X"B1",X"F3",X"A9",X"00",X"A8",X"51",X"30",X"C8",X"D0",
		X"FB",X"60",X"A5",X"31",X"85",X"4E",X"A2",X"01",X"86",X"2F",X"86",X"31",X"CA",X"86",X"4F",X"86",
		X"30",X"20",X"27",X"F9",X"F0",X"0F",X"20",X"E6",X"F7",X"A4",X"36",X"A5",X"52",X"91",X"30",X"C8",
		X"A5",X"53",X"91",X"30",X"C8",X"A5",X"54",X"91",X"30",X"C8",X"A5",X"55",X"91",X"30",X"C8",X"84",
		X"36",X"C0",X"BB",X"90",X"E1",X"A5",X"31",X"85",X"2F",X"A2",X"45",X"86",X"2E",X"A0",X"BB",X"88",
		X"B1",X"30",X"91",X"2E",X"98",X"D0",X"F8",X"A2",X"BB",X"BD",X"00",X"01",X"91",X"30",X"C8",X"E8",
		X"D0",X"F7",X"86",X"50",X"60",X"84",X"36",X"20",X"E6",X"F7",X"A4",X"36",X"A5",X"52",X"91",X"2E",
		X"45",X"4B",X"85",X"4B",X"C8",X"F0",X"ED",X"A5",X"53",X"91",X"2E",X"45",X"4B",X"85",X"4B",X"C8",
		X"A5",X"54",X"91",X"2E",X"45",X"4B",X"85",X"4B",X"C8",X"A5",X"55",X"91",X"2E",X"45",X"4B",X"85",
		X"4B",X"C8",X"D0",X"D1",X"A5",X"85",X"4A",X"C5",X"77",X"F0",X"04",X"C5",X"78",X"D0",X"0D",X"E6",
		X"98",X"A2",X"0F",X"20",X"A5",X"E9",X"CA",X"D0",X"FD",X"20",X"9C",X"E9",X"A2",X"00",X"60",X"50",
		X"60",X"C9",X"20",X"F0",X"03",X"4C",X"CA",X"F6",X"20",X"E9",X"F5",X"85",X"3A",X"20",X"8F",X"F7",
		X"20",X"0A",X"F5",X"A0",X"BB",X"B9",X"00",X"01",X"50",X"FE",X"B8",X"4D",X"01",X"1C",X"D0",X"15",
		X"C8",X"D0",X"F2",X"B1",X"30",X"50",X"FE",X"B8",X"4D",X"01",X"1C",X"D0",X"08",X"C8",X"C0",X"FD",
		X"D0",X"F1",X"4C",X"FE",X"E8",X"A9",X"07",X"4C",X"69",X"F9",X"20",X"10",X"F5",X"4C",X"18",X"F4",
		X"A4",X"34",X"A5",X"53",X"4A",X"4A",X"4A",X"4A",X"AA",X"BD",X"59",X"F7",X"85",X"5A",X"A5",X"52",
		X"29",X"0F",X"AA",X"BD",X"7F",X"F7",X"4A",X"66",X"5A",X"4A",X"66",X"5A",X"85",X"57",X"A5",X"52",
		X"4A",X"4A",X"4A",X"4A",X"AA",X"BD",X"59",X"F7",X"05",X"57",X"91",X"30",X"C8",X"A5",X"53",X"29",
		X"0F",X"AA",X"BD",X"59",X"F7",X"0A",X"85",X"57",X"A5",X"5A",X"69",X"00",X"91",X"30",X"C8",X"A5",
		X"54",X"4A",X"4A",X"4A",X"4A",X"AA",X"BD",X"7F",X"F7",X"4A",X"05",X"57",X"91",X"30",X"C8",X"A5",
		X"54",X"29",X"0F",X"AA",X"BD",X"59",X"F7",X"6A",X"4A",X"4A",X"85",X"5A",X"A5",X"55",X"4A",X"4A",
		X"4A",X"4A",X"AA",X"BD",X"59",X"F7",X"0A",X"26",X"5A",X"0A",X"26",X"5A",X"85",X"57",X"A5",X"5A",
		X"91",X"30",X"C8",X"D0",X"04",X"A5",X"2F",X"85",X"31",X"A5",X"55",X"29",X"0F",X"AA",X"BD",X"7F",
		X"F7",X"05",X"57",X"91",X"30",X"C8",X"84",X"34",X"60",X"50",X"58",X"90",X"98",X"70",X"78",X"B0",
		X"B8",X"48",X"C8",X"D0",X"D8",X"68",X"E8",X"F0",X"A8",X"A5",X"84",X"C9",X"6F",X"B0",X"05",X"20",
		X"25",X"D1",X"90",X"04",X"58",X"4C",X"B7",X"CF",X"A5",X"85",X"4C",X"3A",X"FE",X"34",X"60",X"0A",
		X"0B",X"12",X"13",X"0E",X"0F",X"16",X"17",X"09",X"19",X"1A",X"1B",X"0D",X"1D",X"1E",X"15",X"20",
		X"A6",X"F7",X"85",X"50",X"A5",X"47",X"85",X"52",X"20",X"B9",X"F7",X"A5",X"3A",X"85",X"53",X"84",
		X"54",X"84",X"55",X"4C",X"D0",X"F6",X"A5",X"31",X"85",X"2F",X"A9",X"BB",X"85",X"34",X"A2",X"01",
		X"86",X"31",X"A0",X"00",X"84",X"30",X"84",X"2E",X"60",X"B1",X"2E",X"85",X"53",X"C8",X"B1",X"2E",
		X"85",X"54",X"C8",X"B1",X"2E",X"85",X"55",X"C8",X"F0",X"0E",X"84",X"36",X"20",X"D0",X"F6",X"A4",
		X"36",X"B1",X"2E",X"85",X"52",X"C8",X"D0",X"E1",X"60",X"68",X"C9",X"AF",X"D0",X"06",X"20",X"64",
		X"FB",X"58",X"A9",X"93",X"48",X"60",X"A4",X"34",X"B1",X"30",X"AA",X"29",X"07",X"85",X"57",X"8A",
		X"4A",X"4A",X"4A",X"85",X"56",X"AA",X"C8",X"D0",X"06",X"A5",X"4E",X"85",X"31",X"A4",X"4F",X"B1",
		X"30",X"0A",X"26",X"57",X"0A",X"26",X"57",X"4A",X"4A",X"4A",X"85",X"58",X"BD",X"A0",X"F8",X"A6",
		X"57",X"1D",X"C0",X"F8",X"85",X"52",X"C8",X"B1",X"30",X"6A",X"4A",X"4A",X"4A",X"85",X"59",X"AA",
		X"BD",X"C0",X"F8",X"A6",X"58",X"1D",X"A0",X"F8",X"85",X"53",X"B1",X"30",X"29",X"0F",X"85",X"5A",
		X"C8",X"B1",X"30",X"85",X"5D",X"0A",X"26",X"5A",X"4A",X"4A",X"4A",X"85",X"5B",X"AA",X"BD",X"C0",
		X"F8",X"A6",X"5A",X"1D",X"A0",X"F8",X"85",X"54",X"C8",X"D0",X"06",X"A5",X"4E",X"85",X"31",X"A4",
		X"4F",X"B1",X"30",X"AA",X"46",X"5D",X"6A",X"46",X"5D",X"6A",X"4A",X"4A",X"4A",X"85",X"5C",X"8A",
		X"29",X"1F",X"85",X"5D",X"AA",X"BD",X"C0",X"F8",X"A6",X"5C",X"1D",X"A0",X"F8",X"85",X"55",X"C8",
		X"84",X"34",X"60",X"20",X"E6",X"F7",X"A5",X"52",X"85",X"38",X"A4",X"36",X"4C",X"95",X"F8",X"A5",
		X"54",X"91",X"2E",X"C8",X"A5",X"55",X"91",X"2E",X"C8",X"84",X"36",X"20",X"E6",X"F7",X"A4",X"36",
		X"A5",X"52",X"91",X"2E",X"C8",X"A5",X"53",X"91",X"2E",X"C8",X"D0",X"E3",X"60",X"85",X"55",X"60",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"80",X"00",X"10",X"FF",X"C0",X"40",X"50",
		X"FF",X"FF",X"20",X"30",X"FF",X"F0",X"60",X"70",X"FF",X"90",X"A0",X"B0",X"FF",X"D0",X"E0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"08",X"00",X"01",X"FF",X"0C",X"04",X"05",
		X"FF",X"FF",X"02",X"03",X"FF",X"0F",X"06",X"07",X"FF",X"09",X"0A",X"0B",X"FF",X"0D",X"0E",X"FF",
		X"A2",X"00",X"86",X"36",X"86",X"34",X"86",X"2E",X"86",X"4B",X"E8",X"86",X"4E",X"A2",X"BA",X"86",
		X"4F",X"A6",X"31",X"86",X"2F",X"20",X"01",X"F9",X"A6",X"53",X"86",X"3A",X"A5",X"2F",X"85",X"31",
		X"60",X"20",X"E6",X"F7",X"A5",X"52",X"85",X"38",X"A4",X"36",X"4C",X"57",X"F6",X"20",X"F2",X"F5",
		X"BA",X"BD",X"04",X"01",X"A6",X"3F",X"A0",X"01",X"38",X"E9",X"FB",X"D0",X"E3",X"85",X"50",X"94",
		X"00",X"A6",X"49",X"9A",X"4C",X"BE",X"FA",X"86",X"2E",X"A0",X"BB",X"84",X"36",X"84",X"34",X"4C",
		X"73",X"F8",X"31",X"60",X"A5",X"31",X"85",X"2F",X"A9",X"00",X"85",X"31",X"A9",X"24",X"85",X"34",
		X"A5",X"39",X"85",X"52",X"A5",X"1A",X"85",X"53",X"A5",X"19",X"85",X"54",X"A5",X"18",X"85",X"55",
		X"20",X"D0",X"F6",X"A5",X"17",X"85",X"52",X"A5",X"16",X"85",X"53",X"A9",X"00",X"85",X"54",X"85",
		X"55",X"20",X"D0",X"F6",X"A5",X"2F",X"85",X"31",X"60",X"A4",X"3F",X"99",X"00",X"00",X"A5",X"50",
		X"F0",X"03",X"20",X"F2",X"F5",X"20",X"8F",X"F9",X"A6",X"49",X"9A",X"4C",X"BE",X"F2",X"A9",X"A0",
		X"85",X"20",X"AD",X"00",X"1C",X"09",X"04",X"8D",X"00",X"1C",X"A9",X"19",X"85",X"48",X"60",X"A6",
		X"3E",X"A5",X"20",X"09",X"10",X"85",X"20",X"A9",X"FF",X"85",X"48",X"60",X"AD",X"07",X"1C",X"8D",
		X"05",X"1C",X"AD",X"00",X"1C",X"29",X"10",X"C5",X"1E",X"85",X"1E",X"F0",X"04",X"A9",X"01",X"85",
		X"1C",X"AD",X"FE",X"02",X"F0",X"15",X"C9",X"02",X"D0",X"07",X"A9",X"00",X"8D",X"FE",X"02",X"F0",
		X"0A",X"85",X"4A",X"A9",X"02",X"8D",X"FE",X"02",X"4C",X"2E",X"FA",X"A6",X"3E",X"30",X"07",X"A5",
		X"20",X"A8",X"C9",X"20",X"D0",X"03",X"4C",X"BE",X"FA",X"C6",X"48",X"D0",X"1D",X"98",X"10",X"04",
		X"29",X"7F",X"85",X"20",X"29",X"10",X"F0",X"12",X"AD",X"00",X"1C",X"29",X"FB",X"8D",X"00",X"1C",
		X"A9",X"FF",X"85",X"3E",X"A9",X"00",X"85",X"20",X"F0",X"DC",X"98",X"29",X"40",X"D0",X"03",X"4C",
		X"BE",X"FA",X"6C",X"62",X"00",X"A5",X"4A",X"10",X"05",X"49",X"FF",X"18",X"69",X"01",X"C5",X"64",
		X"B0",X"0A",X"A9",X"3B",X"85",X"62",X"A9",X"FA",X"85",X"63",X"D0",X"12",X"E5",X"5E",X"E5",X"5E",
		X"85",X"61",X"A5",X"5E",X"85",X"60",X"A9",X"7B",X"85",X"62",X"A9",X"FA",X"85",X"63",X"A5",X"4A",
		X"10",X"31",X"E6",X"4A",X"AE",X"00",X"1C",X"CA",X"4C",X"69",X"FA",X"A5",X"4A",X"D0",X"EF",X"A9",
		X"4E",X"85",X"62",X"A9",X"FA",X"85",X"63",X"A9",X"02",X"85",X"60",X"4C",X"BE",X"FA",X"C6",X"60",
		X"D0",X"6C",X"A5",X"20",X"29",X"BF",X"85",X"20",X"A9",X"05",X"85",X"62",X"A9",X"FA",X"85",X"63",
		X"4C",X"BE",X"FA",X"C6",X"4A",X"AE",X"00",X"1C",X"E8",X"8A",X"29",X"03",X"85",X"4B",X"AD",X"00",
		X"1C",X"29",X"FC",X"05",X"4B",X"8D",X"00",X"1C",X"4C",X"BE",X"FA",X"38",X"AD",X"07",X"1C",X"E5",
		X"5F",X"8D",X"05",X"1C",X"C6",X"60",X"D0",X"0C",X"A5",X"5E",X"85",X"60",X"A9",X"97",X"85",X"62",
		X"A9",X"FA",X"85",X"63",X"4C",X"2E",X"FA",X"C6",X"61",X"D0",X"F9",X"A9",X"A5",X"85",X"62",X"A9",
		X"FA",X"85",X"63",X"D0",X"EF",X"AD",X"07",X"1C",X"18",X"65",X"5F",X"8D",X"05",X"1C",X"C6",X"60",
		X"D0",X"E2",X"A9",X"4E",X"85",X"62",X"A9",X"FA",X"85",X"63",X"A9",X"02",X"85",X"60",X"AD",X"0C",
		X"1C",X"29",X"FD",X"8D",X"0C",X"1C",X"60",X"A5",X"51",X"10",X"25",X"20",X"D3",X"FA",X"85",X"51",
		X"4C",X"9C",X"F9",X"A9",X"60",X"85",X"20",X"A9",X"A4",X"85",X"4A",X"A9",X"01",X"85",X"22",X"AD",
		X"00",X"1C",X"29",X"FC",X"8D",X"00",X"1C",X"A9",X"3A",X"8D",X"07",X"1C",X"A9",X"01",X"60",X"AA",
		X"A0",X"00",X"D1",X"32",X"F0",X"05",X"91",X"32",X"4C",X"9C",X"F9",X"A9",X"14",X"8D",X"20",X"06",
		X"AD",X"00",X"1C",X"29",X"10",X"D0",X"05",X"A9",X"08",X"4C",X"DB",X"FD",X"4C",X"3A",X"FC",X"A6",
		X"98",X"30",X"49",X"A4",X"82",X"A1",X"99",X"99",X"3E",X"02",X"B9",X"44",X"02",X"F0",X"0D",X"38",
		X"F5",X"99",X"D0",X"08",X"95",X"99",X"20",X"62",X"D1",X"4C",X"3B",X"FB",X"F6",X"99",X"D0",X"0B",
		X"20",X"74",X"E9",X"20",X"DA",X"D2",X"20",X"2F",X"D1",X"86",X"98",X"A6",X"82",X"AD",X"00",X"18",
		X"29",X"6D",X"85",X"44",X"29",X"61",X"85",X"7A",X"B5",X"F2",X"10",X"A2",X"29",X"08",X"20",X"79",
		X"FF",X"29",X"02",X"F0",X"BA",X"A5",X"7A",X"09",X"0D",X"20",X"DB",X"FF",X"58",X"20",X"AA",X"D3",
		X"78",X"4C",X"3B",X"FB",X"78",X"20",X"D0",X"D6",X"98",X"4A",X"AA",X"A9",X"80",X"20",X"0E",X"D5",
		X"2C",X"A9",X"90",X"48",X"8A",X"0A",X"A8",X"B9",X"06",X"00",X"C5",X"22",X"F0",X"05",X"A9",X"B0",
		X"20",X"A4",X"FB",X"68",X"48",X"95",X"00",X"86",X"3F",X"AD",X"0C",X"1C",X"09",X"0E",X"8D",X"0C",
		X"1C",X"20",X"93",X"F3",X"8A",X"48",X"B5",X"00",X"20",X"AD",X"FB",X"68",X"AA",X"B5",X"00",X"C9",
		X"02",X"68",X"90",X"08",X"20",X"0E",X"D5",X"58",X"20",X"99",X"D5",X"78",X"60",X"BA",X"86",X"49",
		X"29",X"30",X"D0",X"03",X"4C",X"D1",X"F4",X"29",X"20",X"D0",X"03",X"4C",X"75",X"F5",X"4C",X"98",
		X"F6",X"A5",X"98",X"D0",X"03",X"4C",X"C9",X"E9",X"AD",X"00",X"18",X"29",X"04",X"8D",X"00",X"18",
		X"2C",X"00",X"18",X"D0",X"FB",X"48",X"68",X"AD",X"00",X"18",X"0A",X"48",X"68",X"0D",X"00",X"18",
		X"29",X"0F",X"AA",X"A4",X"7A",X"AD",X"00",X"18",X"0A",X"48",X"68",X"0D",X"00",X"18",X"29",X"0F",
		X"1D",X"08",X"FC",X"85",X"85",X"AD",X"00",X"18",X"09",X"02",X"8D",X"00",X"18",X"30",X"C6",X"29",
		X"04",X"D0",X"02",X"84",X"F8",X"A5",X"85",X"60",X"00",X"80",X"20",X"A0",X"40",X"C0",X"60",X"E0",
		X"10",X"90",X"30",X"B0",X"50",X"D0",X"70",X"F0",X"AD",X"0C",X"1C",X"29",X"1F",X"09",X"C0",X"8D",
		X"0C",X"1C",X"A9",X"FF",X"8D",X"03",X"1C",X"60",X"A9",X"FF",X"A2",X"05",X"2C",X"A9",X"55",X"50",
		X"FE",X"B8",X"8D",X"01",X"1C",X"CA",X"D0",X"F7",X"60",X"28",X"8C",X"28",X"06",X"A6",X"3D",X"A5",
		X"39",X"99",X"00",X"03",X"C8",X"C8",X"AD",X"28",X"06",X"99",X"00",X"03",X"C8",X"A5",X"51",X"99",
		X"00",X"03",X"C8",X"B5",X"13",X"99",X"00",X"03",X"C8",X"B5",X"12",X"99",X"00",X"03",X"C8",X"A9",
		X"0F",X"99",X"00",X"03",X"C8",X"99",X"00",X"03",X"C8",X"A9",X"00",X"59",X"FA",X"02",X"59",X"FB",
		X"02",X"59",X"FC",X"02",X"59",X"FD",X"02",X"99",X"F9",X"02",X"EE",X"28",X"06",X"AD",X"28",X"06",
		X"C5",X"43",X"90",X"BB",X"98",X"48",X"E8",X"8A",X"9D",X"00",X"05",X"E8",X"D0",X"FA",X"A9",X"03",
		X"85",X"31",X"20",X"30",X"FE",X"68",X"A8",X"88",X"20",X"E5",X"FD",X"20",X"F5",X"FD",X"A9",X"05",
		X"85",X"31",X"20",X"E9",X"F5",X"85",X"3A",X"20",X"8F",X"F7",X"A5",X"22",X"20",X"4B",X"F2",X"BD",
		X"1A",X"FD",X"AA",X"2C",X"AE",X"26",X"06",X"CA",X"E0",X"04",X"90",X"EE",X"8E",X"26",X"06",X"20",
		X"18",X"FC",X"AA",X"20",X"2D",X"FC",X"86",X"32",X"A5",X"43",X"8D",X"28",X"06",X"A9",X"05",X"85",
		X"31",X"20",X"28",X"FC",X"A2",X"0A",X"A4",X"32",X"50",X"FE",X"B8",X"B9",X"00",X"03",X"8D",X"01",
		X"1C",X"C8",X"CA",X"D0",X"F3",X"A2",X"09",X"20",X"2D",X"FC",X"20",X"28",X"FC",X"A0",X"BB",X"50",
		X"FE",X"B8",X"B9",X"00",X"01",X"8D",X"01",X"1C",X"C8",X"D0",X"F4",X"50",X"FE",X"B8",X"B1",X"30",
		X"8D",X"01",X"1C",X"C8",X"D0",X"F5",X"AE",X"26",X"06",X"20",X"2D",X"FC",X"A5",X"32",X"18",X"69",
		X"0A",X"85",X"32",X"CE",X"28",X"06",X"D0",X"B9",X"F0",X"04",X"08",X"0B",X"10",X"06",X"50",X"FE",
		X"B8",X"50",X"FE",X"B8",X"20",X"00",X"FE",X"A9",X"C8",X"8D",X"23",X"06",X"A9",X"00",X"85",X"30",
		X"A9",X"03",X"85",X"31",X"A5",X"43",X"8D",X"28",X"06",X"20",X"56",X"F5",X"A2",X"0A",X"A0",X"00",
		X"50",X"FE",X"B8",X"AD",X"01",X"1C",X"D1",X"30",X"D0",X"0E",X"C8",X"CA",X"D0",X"F2",X"18",X"A5",
		X"30",X"69",X"0A",X"85",X"30",X"4C",X"62",X"FD",X"CE",X"23",X"06",X"D0",X"CF",X"A9",X"06",X"4C",
		X"D3",X"FD",X"20",X"56",X"F5",X"A0",X"BB",X"50",X"FE",X"B8",X"AD",X"01",X"1C",X"D9",X"00",X"01",
		X"D0",X"E6",X"C8",X"D0",X"F2",X"A2",X"FC",X"50",X"FE",X"B8",X"AD",X"01",X"1C",X"D9",X"00",X"05",
		X"D0",X"D6",X"C8",X"CA",X"D0",X"F1",X"CE",X"28",X"06",X"D0",X"AE",X"E6",X"51",X"A5",X"51",X"C9",
		X"24",X"B0",X"03",X"4C",X"9C",X"F9",X"A9",X"FF",X"85",X"51",X"A9",X"00",X"85",X"50",X"A9",X"01",
		X"4C",X"69",X"F9",X"AD",X"0C",X"1C",X"29",X"1F",X"09",X"C0",X"8D",X"0C",X"1C",X"A9",X"FF",X"8D",
		X"03",X"1C",X"8D",X"01",X"1C",X"A2",X"08",X"A0",X"00",X"50",X"FE",X"B8",X"88",X"D0",X"FA",X"CA",
		X"D0",X"F7",X"60",X"AE",X"21",X"06",X"AC",X"22",X"06",X"50",X"FE",X"B8",X"CA",X"D0",X"FA",X"88",
		X"10",X"F7",X"60",X"CE",X"20",X"06",X"F0",X"03",X"4C",X"B4",X"FC",X"A0",X"FF",X"84",X"51",X"C8",
		X"84",X"50",X"4C",X"69",X"F9",X"B9",X"00",X"03",X"99",X"45",X"03",X"88",X"D0",X"F7",X"AD",X"00",
		X"03",X"8D",X"45",X"03",X"60",X"A0",X"44",X"B9",X"BB",X"01",X"91",X"30",X"88",X"10",X"F8",X"60",
		X"AD",X"0C",X"1C",X"09",X"E0",X"8D",X"0C",X"1C",X"A9",X"00",X"8D",X"03",X"1C",X"60",X"AD",X"0C",
		X"1C",X"29",X"1F",X"09",X"C0",X"8D",X"0C",X"1C",X"A9",X"FF",X"8D",X"03",X"1C",X"A9",X"55",X"8D",
		X"01",X"1C",X"A2",X"08",X"A0",X"00",X"50",X"FE",X"B8",X"88",X"D0",X"FA",X"CA",X"D0",X"F7",X"60",
		X"20",X"A6",X"F7",X"20",X"D1",X"F7",X"4C",X"D0",X"F6",X"BB",X"20",X"F1",X"CF",X"D0",X"27",X"20",
		X"B7",X"DF",X"D0",X"05",X"58",X"20",X"7B",X"CF",X"78",X"29",X"07",X"AA",X"B5",X"00",X"10",X"03",
		X"20",X"73",X"FB",X"58",X"20",X"1E",X"F1",X"78",X"20",X"A9",X"D1",X"A6",X"F9",X"20",X"71",X"FB",
		X"A6",X"F9",X"A9",X"A0",X"95",X"00",X"60",X"48",X"8A",X"48",X"98",X"48",X"AD",X"0D",X"18",X"29",
		X"02",X"F0",X"03",X"20",X"53",X"E8",X"AD",X"0D",X"1C",X"0A",X"10",X"03",X"20",X"B0",X"F2",X"68",
		X"A8",X"68",X"AA",X"68",X"40",X"12",X"04",X"04",X"90",X"56",X"49",X"44",X"4D",X"42",X"55",X"50",
		X"26",X"43",X"52",X"53",X"4E",X"84",X"05",X"C1",X"F8",X"1B",X"5C",X"07",X"A3",X"F0",X"88",X"23",
		X"0D",X"ED",X"D0",X"C8",X"CA",X"CC",X"CB",X"E2",X"E7",X"C8",X"CA",X"C8",X"EE",X"51",X"DD",X"1C",
		X"9E",X"1C",X"52",X"57",X"41",X"4D",X"44",X"53",X"50",X"55",X"4C",X"44",X"53",X"50",X"55",X"52",
		X"45",X"45",X"52",X"53",X"45",X"4C",X"51",X"47",X"52",X"4C",X"08",X"00",X"00",X"3F",X"7F",X"BF",
		X"FF",X"11",X"12",X"13",X"15",X"41",X"04",X"24",X"1F",X"19",X"12",X"01",X"FF",X"FF",X"01",X"00",
		X"03",X"04",X"05",X"06",X"07",X"07",X"BB",X"6C",X"65",X"00",X"8D",X"00",X"1C",X"8D",X"02",X"1C",
		X"4C",X"7D",X"EA",X"8A",X"A2",X"05",X"CA",X"D0",X"FD",X"AA",X"60",X"20",X"AE",X"E9",X"4C",X"9C",
		X"E9",X"AD",X"02",X"02",X"C9",X"2D",X"F0",X"05",X"38",X"E9",X"2B",X"D0",X"DA",X"85",X"23",X"60",
		X"8E",X"03",X"18",X"A9",X"02",X"8D",X"00",X"18",X"A9",X"1A",X"8D",X"02",X"18",X"4C",X"A7",X"EA",
		X"AD",X"00",X"18",X"29",X"01",X"D0",X"F9",X"A9",X"01",X"8D",X"05",X"18",X"60",X"A5",X"31",X"48",
		X"20",X"6D",X"E9",X"A9",X"04",X"48",X"A0",X"01",X"B1",X"30",X"85",X"81",X"AA",X"88",X"B1",X"30",
		X"85",X"80",X"D0",X"0C",X"68",X"18",X"E5",X"81",X"E8",X"86",X"30",X"F0",X"02",X"C6",X"31",X"48",
		X"68",X"A8",X"20",X"8D",X"FF",X"A5",X"80",X"F0",X"07",X"20",X"64",X"FB",X"A9",X"02",X"D0",X"D5",
		X"85",X"30",X"68",X"85",X"31",X"20",X"6E",X"FF",X"20",X"6E",X"FF",X"20",X"AE",X"E9",X"A2",X"14",
		X"CA",X"D0",X"FD",X"4C",X"B7",X"E9",X"4C",X"5B",X"E8",X"D0",X"06",X"A5",X"7A",X"09",X"03",X"85",
		X"44",X"BD",X"3E",X"02",X"A6",X"7A",X"A0",X"FF",X"8E",X"00",X"18",X"D0",X"18",X"AD",X"00",X"18",
		X"29",X"60",X"85",X"7A",X"09",X"0D",X"85",X"44",X"20",X"A5",X"E9",X"49",X"0D",X"8D",X"00",X"18",
		X"20",X"F3",X"FE",X"B1",X"30",X"AA",X"4A",X"4A",X"4A",X"4A",X"85",X"4B",X"8A",X"29",X"0F",X"AA",
		X"BD",X"1D",X"EA",X"A6",X"7A",X"8E",X"00",X"18",X"EC",X"00",X"18",X"F0",X"FB",X"8D",X"00",X"18",
		X"0A",X"29",X"0F",X"EA",X"8D",X"00",X"18",X"A6",X"4B",X"BD",X"1D",X"EA",X"8D",X"00",X"18",X"0A",
		X"29",X"0F",X"C8",X"8D",X"00",X"18",X"D0",X"CB",X"EA",X"A5",X"44",X"8D",X"00",X"18",X"CD",X"00",
		X"18",X"90",X"93",X"D0",X"F9",X"60",X"C6",X"C8",X"8F",X"F9",X"5F",X"CD",X"97",X"CD",X"00",X"05",
		X"03",X"05",X"06",X"05",X"09",X"05",X"0C",X"05",X"0F",X"05",X"01",X"FF",X"A0",X"EA",X"67",X"FE");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
