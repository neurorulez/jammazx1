library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_pgme is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_pgme is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"D2",X"74",X"D3",X"12",X"D2",X"CC",X"D3",X"30",X"D2",X"33",X"D2",X"36",X"CF",X"D7",X"D1",X"36",
		X"CF",X"26",X"D2",X"36",X"CF",X"EE",X"D3",X"36",X"CF",X"36",X"CF",X"21",X"D4",X"36",X"CF",X"36",
		X"CF",X"36",X"CF",X"4E",X"D2",X"36",X"CF",X"36",X"CF",X"90",X"D4",X"BC",X"D4",X"F1",X"D3",X"36",
		X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",
		X"CF",X"36",X"CF",X"36",X"CF",X"65",X"D3",X"50",X"D4",X"33",X"D4",X"24",X"D4",X"2E",X"D1",X"48",
		X"D1",X"09",X"D4",X"36",X"CF",X"D7",X"D1",X"3C",X"D4",X"3C",X"D4",X"36",X"CF",X"36",X"CF",X"36",
		X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"90",X"D4",X"BC",X"D4",X"36",
		X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"90",X"D4",X"BC",
		X"D4",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"0A",X"D3",X"36",X"CF",X"36",X"CF",X"90",X"D4",X"BC",
		X"D4",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",
		X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",
		X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"36",X"CF",X"90",X"D4",X"BC",X"D4",X"36",X"CF",X"36",
		X"CF",X"36",X"CF",X"90",X"D4",X"BC",X"D4",X"BC",X"D4",X"8A",X"A8",X"4C",X"13",X"D2",X"4C",X"37",
		X"CF",X"BD",X"0A",X"02",X"85",X"59",X"BD",X"0C",X"02",X"85",X"5B",X"A9",X"07",X"85",X"5D",X"20",
		X"03",X"D5",X"B0",X"09",X"A9",X"00",X"85",X"5D",X"20",X"1F",X"D5",X"B0",X"10",X"A9",X"03",X"99",
		X"00",X"02",X"20",X"78",X"D3",X"A9",X"00",X"20",X"46",X"C8",X"4C",X"37",X"CF",X"A9",X"00",X"9D",
		X"00",X"21",X"9D",X"06",X"21",X"A9",X"0B",X"9D",X"01",X"02",X"A9",X"1F",X"9D",X"0D",X"02",X"A9",
		X"25",X"84",X"19",X"A9",X"00",X"9D",X"00",X"02",X"A8",X"20",X"1B",X"CA",X"A4",X"19",X"20",X"2A",
		X"BD",X"A9",X"03",X"99",X"00",X"02",X"4C",X"37",X"CF",X"4C",X"37",X"CF",X"4C",X"37",X"CF",X"B9",
		X"01",X"02",X"29",X"F0",X"09",X"0A",X"99",X"01",X"02",X"A9",X"01",X"99",X"0D",X"02",X"A9",X"03",
		X"9D",X"00",X"02",X"20",X"2A",X"BD",X"4C",X"37",X"CF",X"A9",X"03",X"9D",X"00",X"02",X"EE",X"03",
		X"03",X"AD",X"03",X"03",X"C9",X"0B",X"D0",X"03",X"4C",X"65",X"D1",X"98",X"AA",X"A9",X"09",X"20",
		X"46",X"C8",X"4C",X"37",X"CF",X"A6",X"41",X"86",X"19",X"A9",X"00",X"9D",X"01",X"02",X"A9",X"00",
		X"85",X"59",X"A9",X"50",X"85",X"5A",X"A9",X"00",X"85",X"5B",X"20",X"80",X"D1",X"4C",X"37",X"CF",
		X"A9",X"60",X"9D",X"01",X"21",X"A9",X"00",X"9D",X"00",X"21",X"9D",X"06",X"21",X"A5",X"5B",X"24",
		X"EF",X"30",X"20",X"F8",X"18",X"6D",X"43",X"04",X"8D",X"43",X"04",X"A5",X"5A",X"6D",X"42",X"04",
		X"8D",X"42",X"04",X"A5",X"59",X"6D",X"41",X"04",X"8D",X"41",X"04",X"D8",X"A0",X"00",X"A9",X"00",
		X"20",X"1B",X"CA",X"20",X"AD",X"C8",X"60",X"98",X"AA",X"A9",X"00",X"20",X"46",X"C8",X"4C",X"37",
		X"CF",X"A9",X"01",X"99",X"00",X"02",X"A9",X"14",X"99",X"0D",X"02",X"A0",X"00",X"A9",X"25",X"20",
		X"1B",X"CA",X"20",X"2A",X"BD",X"4C",X"37",X"CF",X"A5",X"73",X"D0",X"F9",X"B9",X"00",X"02",X"29",
		X"03",X"D0",X"F2",X"A9",X"01",X"99",X"00",X"02",X"A9",X"00",X"99",X"03",X"02",X"A9",X"01",X"99",
		X"0D",X"02",X"99",X"02",X"02",X"A9",X"00",X"99",X"00",X"21",X"99",X"06",X"21",X"AD",X"64",X"56",
		X"99",X"04",X"21",X"AD",X"65",X"56",X"99",X"05",X"21",X"A0",X"05",X"A9",X"00",X"20",X"1B",X"CA",
		X"4C",X"37",X"CF",X"A5",X"6C",X"D0",X"0D",X"A5",X"73",X"D0",X"09",X"84",X"6C",X"20",X"0E",X"BE",
		X"20",X"52",X"BD",X"60",X"4C",X"37",X"CF",X"B9",X"00",X"02",X"29",X"03",X"D0",X"F6",X"4C",X"13",
		X"D2",X"4C",X"13",X"D2",X"20",X"9B",X"D3",X"98",X"AA",X"B9",X"0D",X"02",X"29",X"18",X"4A",X"4A",
		X"4A",X"A8",X"B9",X"4B",X"D2",X"20",X"46",X"C8",X"4C",X"37",X"CF",X"01",X"03",X"09",X"13",X"AD",
		X"0A",X"60",X"10",X"03",X"4C",X"AC",X"D2",X"A9",X"08",X"9D",X"00",X"02",X"20",X"3E",X"BD",X"A9",
		X"14",X"9D",X"0D",X"02",X"B9",X"09",X"02",X"9D",X"09",X"02",X"B9",X"0A",X"02",X"9D",X"0A",X"02",
		X"B9",X"0B",X"02",X"9D",X"0B",X"02",X"B9",X"0C",X"02",X"9D",X"0C",X"02",X"B9",X"01",X"02",X"29",
		X"F0",X"09",X"03",X"99",X"01",X"02",X"99",X"02",X"02",X"A9",X"03",X"99",X"0F",X"02",X"A9",X"00",
		X"99",X"00",X"02",X"A9",X"1F",X"99",X"0D",X"02",X"A9",X"00",X"99",X"02",X"21",X"A9",X"73",X"99",
		X"03",X"21",X"84",X"40",X"A9",X"00",X"99",X"00",X"02",X"4C",X"37",X"CF",X"86",X"19",X"98",X"AA",
		X"A4",X"19",X"A9",X"01",X"25",X"9A",X"F0",X"50",X"20",X"3E",X"BD",X"B9",X"00",X"02",X"09",X"08",
		X"99",X"00",X"02",X"A9",X"14",X"99",X"0D",X"02",X"BD",X"09",X"02",X"99",X"09",X"02",X"BD",X"0A",
		X"02",X"99",X"0A",X"02",X"BD",X"0B",X"02",X"99",X"0B",X"02",X"BD",X"0C",X"02",X"99",X"0C",X"02",
		X"BD",X"01",X"02",X"29",X"F0",X"09",X"03",X"9D",X"01",X"02",X"A9",X"03",X"9D",X"0F",X"02",X"A9",
		X"00",X"9D",X"02",X"02",X"9D",X"00",X"02",X"A9",X"1F",X"9D",X"0D",X"02",X"A9",X"00",X"9D",X"02",
		X"21",X"A9",X"73",X"9D",X"03",X"21",X"86",X"40",X"4C",X"37",X"CF",X"A9",X"03",X"99",X"00",X"02",
		X"20",X"36",X"BD",X"4C",X"37",X"CF",X"B9",X"00",X"02",X"29",X"F7",X"99",X"00",X"02",X"84",X"40",
		X"B9",X"06",X"02",X"48",X"BD",X"07",X"02",X"99",X"07",X"02",X"BD",X"08",X"02",X"99",X"08",X"02",
		X"BD",X"06",X"02",X"99",X"06",X"02",X"20",X"EE",X"C3",X"A6",X"40",X"68",X"9D",X"06",X"02",X"4C",
		X"37",X"CF",X"A5",X"73",X"F0",X"1D",X"A9",X"00",X"85",X"73",X"8D",X"03",X"03",X"8D",X"01",X"03",
		X"24",X"EF",X"30",X"0F",X"A9",X"E4",X"8D",X"02",X"01",X"8D",X"03",X"01",X"AD",X"06",X"02",X"49",
		X"FF",X"85",X"72",X"4C",X"37",X"CF",X"A9",X"03",X"9D",X"00",X"02",X"98",X"AA",X"A9",X"22",X"20",
		X"46",X"C8",X"4C",X"37",X"CF",X"4C",X"13",X"D2",X"AD",X"04",X"03",X"F0",X"1D",X"86",X"19",X"86",
		X"1B",X"84",X"1C",X"85",X"1D",X"AA",X"BD",X"04",X"03",X"A8",X"B9",X"02",X"02",X"C5",X"19",X"F0",
		X"14",X"CA",X"C6",X"1D",X"D0",X"F0",X"A6",X"1B",X"A4",X"1C",X"60",X"AD",X"04",X"03",X"F0",X"FA",
		X"84",X"19",X"4C",X"7F",X"D3",X"A9",X"00",X"99",X"02",X"02",X"68",X"68",X"A6",X"19",X"AD",X"D3",
		X"03",X"0A",X"69",X"17",X"C9",X"20",X"90",X"02",X"A9",X"1F",X"20",X"46",X"C8",X"EE",X"D3",X"03",
		X"4C",X"37",X"CF",X"A5",X"73",X"F0",X"03",X"4C",X"37",X"CF",X"4C",X"13",X"D2",X"4C",X"13",X"D2",
		X"AD",X"0A",X"60",X"29",X"30",X"18",X"7D",X"0E",X"02",X"29",X"3F",X"9D",X"0E",X"02",X"4C",X"37",
		X"CF",X"BD",X"00",X"02",X"29",X"F7",X"9D",X"00",X"02",X"20",X"DE",X"C3",X"4C",X"37",X"CF",X"4C",
		X"D1",X"D0",X"AD",X"0A",X"60",X"29",X"87",X"10",X"02",X"09",X"F8",X"18",X"79",X"06",X"02",X"29",
		X"3F",X"99",X"06",X"02",X"20",X"2A",X"BD",X"4C",X"37",X"CF",X"AD",X"0A",X"60",X"29",X"87",X"10",
		X"02",X"09",X"F8",X"18",X"7D",X"06",X"02",X"29",X"3F",X"9D",X"06",X"02",X"20",X"2A",X"BD",X"4C",
		X"37",X"CF",X"4C",X"37",X"CF",X"A9",X"03",X"9D",X"00",X"02",X"98",X"AA",X"A9",X"20",X"20",X"46",
		X"C8",X"4C",X"37",X"CF",X"98",X"48",X"8A",X"A8",X"68",X"AA",X"4C",X"D1",X"D0",X"B9",X"00",X"02",
		X"29",X"01",X"D0",X"39",X"B9",X"05",X"02",X"18",X"69",X"01",X"C9",X"10",X"B0",X"03",X"99",X"05",
		X"02",X"A9",X"03",X"9D",X"00",X"02",X"B9",X"06",X"02",X"48",X"BD",X"07",X"02",X"99",X"07",X"02",
		X"BD",X"08",X"02",X"99",X"08",X"02",X"BD",X"06",X"02",X"99",X"06",X"02",X"84",X"40",X"20",X"EE",
		X"C3",X"A6",X"40",X"68",X"9D",X"06",X"02",X"20",X"2A",X"BD",X"4C",X"37",X"CF",X"A9",X"03",X"9D",
		X"00",X"02",X"A9",X"00",X"99",X"01",X"02",X"98",X"AA",X"A9",X"20",X"20",X"46",X"C8",X"4C",X"37",
		X"CF",X"8A",X"D9",X"02",X"02",X"D0",X"F7",X"BD",X"00",X"02",X"29",X"03",X"C9",X"02",X"B0",X"1A",
		X"A9",X"03",X"9D",X"00",X"02",X"AD",X"3F",X"04",X"0A",X"99",X"0D",X"02",X"A9",X"00",X"8D",X"D3",
		X"03",X"99",X"02",X"02",X"99",X"05",X"02",X"20",X"36",X"BD",X"4C",X"37",X"CF",X"BD",X"00",X"02",
		X"29",X"03",X"C9",X"02",X"B0",X"3A",X"BD",X"01",X"02",X"29",X"0F",X"C9",X"05",X"D0",X"09",X"A5",
		X"79",X"C9",X"1E",X"B0",X"03",X"4C",X"37",X"CF",X"BD",X"01",X"02",X"29",X"F0",X"09",X"08",X"9D",
		X"01",X"02",X"A9",X"71",X"9D",X"03",X"21",X"9D",X"0B",X"21",X"A9",X"FF",X"9D",X"02",X"02",X"9D",
		X"04",X"02",X"A9",X"00",X"9D",X"0A",X"21",X"9D",X"00",X"02",X"9D",X"0D",X"02",X"20",X"26",X"BD",
		X"4C",X"37",X"CF",X"A5",X"59",X"10",X"06",X"49",X"FF",X"85",X"59",X"E6",X"59",X"A5",X"5B",X"10",
		X"06",X"49",X"FF",X"85",X"5B",X"E6",X"5B",X"A5",X"59",X"85",X"5A",X"A5",X"5B",X"85",X"5C",X"84",
		X"19",X"A5",X"5D",X"0A",X"0A",X"65",X"5D",X"65",X"5D",X"A8",X"B9",X"6F",X"BF",X"C5",X"59",X"90",
		X"21",X"B9",X"71",X"BF",X"C5",X"5B",X"90",X"1A",X"A5",X"59",X"4A",X"18",X"65",X"5B",X"D9",X"6F",
		X"BF",X"B0",X"0F",X"A5",X"59",X"0A",X"18",X"65",X"5B",X"D9",X"73",X"BF",X"B0",X"04",X"18",X"A4",
		X"19",X"60",X"38",X"A4",X"19",X"60",X"27",X"2C",X"30",X"34",X"39",X"00",X"07",X"0C",X"10",X"14",
		X"19",X"20",X"61",X"00",X"A2",X"02",X"AD",X"00",X"78",X"E0",X"01",X"F0",X"03",X"B0",X"02",X"4A",
		X"4A",X"4A",X"B5",X"91",X"29",X"1F",X"B0",X"37",X"F0",X"10",X"C9",X"1B",X"B0",X"0A",X"A8",X"A5",
		X"94",X"29",X"07",X"C9",X"07",X"98",X"90",X"02",X"E9",X"01",X"95",X"91",X"AD",X"00",X"78",X"29",
		X"08",X"D0",X"04",X"A9",X"F0",X"85",X"96",X"A5",X"96",X"F0",X"08",X"C6",X"96",X"A9",X"00",X"95",
		X"91",X"95",X"8E",X"18",X"B5",X"8E",X"F0",X"23",X"D6",X"8E",X"D0",X"1F",X"38",X"B0",X"1C",X"C9",
		X"1B",X"B0",X"09",X"B5",X"91",X"69",X"20",X"90",X"D1",X"F0",X"01",X"18",X"A9",X"1F",X"B0",X"CA",
		X"95",X"91",X"B5",X"8E",X"F0",X"01",X"38",X"A9",X"78",X"95",X"8E",X"90",X"2A",X"A9",X"00",X"E0",
		X"01",X"90",X"16",X"F0",X"0C",X"A5",X"8C",X"29",X"0C",X"4A",X"4A",X"F0",X"0C",X"69",X"02",X"D0",
		X"08",X"A5",X"8C",X"29",X"10",X"F0",X"02",X"A9",X"01",X"38",X"48",X"65",X"F5",X"85",X"F5",X"68",
		X"38",X"65",X"95",X"85",X"95",X"F6",X"89",X"CA",X"30",X"03",X"4C",X"66",X"D5",X"A5",X"8C",X"4A",
		X"4A",X"4A",X"4A",X"4A",X"A8",X"A5",X"F5",X"38",X"F9",X"19",X"D6",X"30",X"14",X"85",X"F5",X"E6",
		X"F4",X"C0",X"03",X"D0",X"0C",X"E6",X"F4",X"D0",X"08",X"7F",X"02",X"04",X"04",X"05",X"03",X"7F",
		X"7F",X"A5",X"8C",X"29",X"03",X"A8",X"F0",X"1A",X"4A",X"69",X"00",X"49",X"FF",X"38",X"65",X"95",
		X"B0",X"08",X"65",X"F4",X"30",X"0E",X"85",X"F4",X"A9",X"00",X"C0",X"02",X"B0",X"02",X"E6",X"8D",
		X"E6",X"8D",X"85",X"95",X"A5",X"94",X"4A",X"B0",X"27",X"A0",X"00",X"A2",X"02",X"B5",X"89",X"F0",
		X"09",X"C9",X"10",X"90",X"05",X"69",X"EF",X"C8",X"95",X"89",X"CA",X"10",X"F0",X"98",X"D0",X"10",
		X"A2",X"02",X"B5",X"89",X"F0",X"07",X"18",X"69",X"EF",X"95",X"89",X"30",X"03",X"CA",X"10",X"F2",
		X"60",X"00",X"02",X"03",X"18",X"19",X"1C",X"1D",X"20",X"7A",X"00",X"10",X"03",X"76",X"00",X"7C",
		X"00",X"A9",X"04",X"D0",X"06",X"A9",X"03",X"D0",X"02",X"A9",X"07",X"A0",X"FF",X"D0",X"08",X"A9",
		X"02",X"D0",X"02",X"A9",X"0D",X"A0",X"00",X"8C",X"2A",X"01",X"48",X"0D",X"2B",X"01",X"8D",X"2B",
		X"01",X"68",X"0D",X"2C",X"01",X"8D",X"2C",X"01",X"60",X"A9",X"0F",X"8D",X"2B",X"01",X"A9",X"00",
		X"8D",X"2C",X"01",X"AD",X"2E",X"01",X"D0",X"4B",X"AD",X"2B",X"01",X"F0",X"46",X"A2",X"00",X"8E",
		X"2F",X"01",X"8E",X"33",X"01",X"8E",X"32",X"01",X"A2",X"08",X"38",X"6E",X"32",X"01",X"0A",X"CA",
		X"90",X"F9",X"A0",X"80",X"AD",X"32",X"01",X"2D",X"2C",X"01",X"D0",X"02",X"A0",X"20",X"8C",X"2E",
		X"01",X"AD",X"32",X"01",X"4D",X"2B",X"01",X"8D",X"2B",X"01",X"8A",X"0A",X"AA",X"BD",X"71",X"D6",
		X"8D",X"30",X"01",X"BD",X"72",X"D6",X"8D",X"31",X"01",X"BD",X"79",X"D6",X"85",X"97",X"BD",X"7A",
		X"D6",X"85",X"98",X"A0",X"00",X"8C",X"00",X"89",X"AD",X"2E",X"01",X"D0",X"01",X"60",X"AC",X"2F",
		X"01",X"AE",X"30",X"01",X"0A",X"90",X"0D",X"9D",X"40",X"89",X"A9",X"40",X"8D",X"2E",X"01",X"A0",
		X"0E",X"4C",X"98",X"D7",X"10",X"25",X"A9",X"80",X"8D",X"2E",X"01",X"AD",X"2A",X"01",X"F0",X"04",
		X"A9",X"00",X"91",X"97",X"B1",X"97",X"EC",X"31",X"01",X"90",X"08",X"A9",X"00",X"8D",X"2E",X"01",
		X"AD",X"33",X"01",X"9D",X"40",X"89",X"A0",X"0C",X"4C",X"8B",X"D7",X"A9",X"08",X"8D",X"00",X"89",
		X"9D",X"40",X"89",X"A9",X"09",X"8D",X"00",X"89",X"EA",X"A9",X"08",X"8D",X"00",X"89",X"EC",X"31",
		X"01",X"AD",X"00",X"70",X"90",X"21",X"4D",X"33",X"01",X"F0",X"14",X"A9",X"00",X"AC",X"2F",X"01",
		X"88",X"91",X"97",X"88",X"10",X"FB",X"AD",X"32",X"01",X"0D",X"2D",X"01",X"8D",X"2D",X"01",X"A9",
		X"00",X"8D",X"2E",X"01",X"4C",X"89",X"D7",X"91",X"97",X"A0",X"00",X"18",X"6D",X"33",X"01",X"8D",
		X"33",X"01",X"EE",X"2F",X"01",X"EE",X"30",X"01",X"8C",X"00",X"89",X"98",X"D0",X"03",X"4C",X"B3",
		X"D6",X"60",X"A9",X"C0",X"D0",X"02",X"A9",X"20",X"A0",X"00",X"91",X"11",X"4C",X"54",X"D8",X"90",
		X"04",X"29",X"0F",X"F0",X"05",X"29",X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",
		X"C4",X"5D",X"91",X"11",X"BD",X"C5",X"5D",X"C8",X"91",X"11",X"20",X"05",X"D8",X"28",X"60",X"38",
		X"E9",X"20",X"4A",X"29",X"1F",X"09",X"E0",X"A0",X"01",X"91",X"11",X"88",X"8A",X"6A",X"91",X"11",
		X"C8",X"D0",X"22",X"38",X"E9",X"20",X"4A",X"29",X"1F",X"09",X"A0",X"D0",X"EA",X"A4",X"0C",X"A2",
		X"60",X"98",X"4C",X"FD",X"D7",X"A2",X"60",X"D0",X"F8",X"A9",X"40",X"A2",X"80",X"A0",X"00",X"91",
		X"11",X"C8",X"8A",X"91",X"11",X"98",X"38",X"65",X"11",X"85",X"11",X"90",X"02",X"E6",X"12",X"60",
		X"A0",X"00",X"09",X"70",X"AA",X"98",X"4C",X"FD",X"D7",X"A0",X"00",X"84",X"0C",X"A0",X"00",X"0A",
		X"90",X"01",X"88",X"84",X"A0",X"0A",X"26",X"A0",X"85",X"9F",X"8A",X"0A",X"A0",X"00",X"90",X"01",
		X"88",X"84",X"A2",X"0A",X"26",X"A2",X"85",X"A1",X"A2",X"9F",X"A0",X"00",X"B5",X"02",X"91",X"11",
		X"B5",X"03",X"29",X"1F",X"C8",X"91",X"11",X"B5",X"00",X"C8",X"91",X"11",X"B5",X"01",X"45",X"0C",
		X"29",X"1F",X"45",X"0C",X"C8",X"91",X"11",X"D0",X"AC",X"A5",X"0C",X"A0",X"00",X"91",X"11",X"C8",
		X"8A",X"09",X"60",X"91",X"11",X"20",X"05",X"D8",X"60",X"00",X"00",X"D0",X"1F",X"4E",X"BE",X"4E",
		X"BE",X"4E",X"BE",X"4E",X"BE",X"4E",X"BE",X"00",X"C0",X"48",X"A5",X"74",X"85",X"4C",X"A5",X"75",
		X"85",X"4D",X"A9",X"04",X"CA",X"30",X"06",X"18",X"69",X"06",X"4C",X"84",X"D8",X"A8",X"68",X"38",
		X"E9",X"02",X"F0",X"0D",X"AA",X"98",X"18",X"69",X"4E",X"90",X"02",X"E6",X"4D",X"CA",X"D0",X"F6",
		X"A8",X"60",X"A9",X"06",X"85",X"19",X"A9",X"A4",X"AA",X"A9",X"5C",X"20",X"E3",X"D7",X"C6",X"19",
		X"D0",X"F4",X"60",X"A8",X"A1",X"B0",X"A1",X"B8",X"A1",X"C0",X"A1",X"C8",X"A1",X"D0",X"A1",X"D8",
		X"A1",X"E0",X"A1",X"E8",X"A1",X"F0",X"A1",X"F8",X"A1",X"A0",X"00",X"A9",X"80",X"91",X"11",X"C8",
		X"A9",X"80",X"91",X"11",X"20",X"05",X"D8",X"A9",X"00",X"85",X"0D",X"85",X"0F",X"85",X"0E",X"85",
		X"10",X"60",X"A9",X"FF",X"4C",X"E9",X"D8",X"A9",X"00",X"48",X"A2",X"00",X"38",X"B5",X"08",X"A8",
		X"F5",X"0D",X"95",X"08",X"98",X"95",X"0D",X"E8",X"B5",X"08",X"A8",X"F5",X"0D",X"95",X"08",X"98",
		X"95",X"0D",X"E8",X"E0",X"02",X"F0",X"E5",X"68",X"D0",X"45",X"A0",X"00",X"A2",X"03",X"98",X"15",
		X"08",X"A8",X"CA",X"10",X"F9",X"98",X"F0",X"37",X"A2",X"02",X"B5",X"09",X"10",X"0F",X"49",X"FF",
		X"D0",X"2D",X"B5",X"08",X"49",X"FF",X"18",X"69",X"01",X"B0",X"24",X"90",X"02",X"B5",X"08",X"29",
		X"1F",X"D0",X"1C",X"B5",X"08",X"29",X"1F",X"95",X"08",X"CA",X"CA",X"10",X"DD",X"A5",X"0C",X"05",
		X"08",X"A0",X"00",X"91",X"11",X"C8",X"A5",X"0A",X"09",X"40",X"91",X"11",X"4C",X"05",X"D8",X"20",
		X"56",X"D9",X"20",X"05",X"D8",X"60",X"A0",X"00",X"A5",X"0A",X"91",X"11",X"C8",X"A5",X"0B",X"29",
		X"1F",X"91",X"11",X"C8",X"A5",X"08",X"91",X"11",X"C8",X"A5",X"09",X"29",X"1F",X"05",X"0C",X"91",
		X"11",X"60",X"A5",X"AA",X"85",X"11",X"A5",X"AB",X"85",X"12",X"24",X"EF",X"10",X"3C",X"AD",X"20",
		X"04",X"C9",X"01",X"D0",X"0F",X"A5",X"F7",X"C9",X"08",X"B0",X"09",X"4A",X"AA",X"BD",X"5C",X"DA",
		X"AA",X"20",X"B7",X"DC",X"A9",X"EC",X"85",X"59",X"A9",X"60",X"85",X"5B",X"AD",X"75",X"CB",X"85",
		X"63",X"A9",X"40",X"85",X"5A",X"AD",X"77",X"CB",X"85",X"5C",X"A2",X"00",X"86",X"19",X"A0",X"00",
		X"20",X"3B",X"CD",X"88",X"20",X"05",X"D8",X"4C",X"15",X"DA",X"AD",X"C8",X"04",X"F0",X"0E",X"AD",
		X"C9",X"04",X"F0",X"09",X"AD",X"40",X"04",X"8D",X"AA",X"04",X"4C",X"D3",X"D9",X"AD",X"40",X"04",
		X"8D",X"75",X"04",X"AD",X"45",X"04",X"F0",X"3A",X"A2",X"34",X"20",X"B7",X"DC",X"AD",X"47",X"04",
		X"85",X"1E",X"A9",X"00",X"F8",X"18",X"6D",X"45",X"04",X"C6",X"1E",X"10",X"F8",X"D8",X"85",X"1B",
		X"4A",X"4A",X"4A",X"4A",X"F0",X"03",X"20",X"AF",X"D7",X"A5",X"1B",X"20",X"AF",X"D7",X"A9",X"00",
		X"20",X"AF",X"D7",X"A9",X"00",X"20",X"AF",X"D7",X"A9",X"00",X"20",X"AF",X"D7",X"A9",X"00",X"20",
		X"AF",X"D7",X"4C",X"34",X"DA",X"20",X"6F",X"DE",X"A2",X"2A",X"20",X"B7",X"DC",X"A5",X"8C",X"29",
		X"03",X"F0",X"0C",X"A5",X"8D",X"D0",X"08",X"A2",X"20",X"20",X"B7",X"DC",X"4C",X"34",X"DA",X"A2",
		X"06",X"20",X"B7",X"DC",X"24",X"EF",X"30",X"1D",X"A2",X"1A",X"20",X"B7",X"DC",X"AD",X"5D",X"04",
		X"18",X"69",X"01",X"20",X"A1",X"DC",X"48",X"4A",X"4A",X"4A",X"4A",X"38",X"20",X"AF",X"D7",X"68",
		X"29",X"0F",X"20",X"AF",X"D7",X"20",X"A2",X"D7",X"20",X"87",X"CA",X"60",X"58",X"5A",X"5C",X"5E",
		X"18",X"F0",X"05",X"C6",X"1C",X"4C",X"AF",X"D7",X"24",X"1C",X"30",X"01",X"38",X"4C",X"AF",X"D7",
		X"A5",X"AA",X"85",X"11",X"A5",X"AB",X"85",X"12",X"A9",X"00",X"A2",X"28",X"20",X"1D",X"D8",X"A9",
		X"00",X"20",X"10",X"D8",X"AD",X"5D",X"04",X"29",X"78",X"4A",X"4A",X"C9",X"0A",X"90",X"02",X"A9",
		X"08",X"AA",X"A0",X"00",X"BD",X"66",X"56",X"91",X"11",X"C8",X"BD",X"67",X"56",X"91",X"11",X"E6",
		X"11",X"E6",X"11",X"20",X"F9",X"D7",X"A9",X"01",X"20",X"10",X"D8",X"A9",X"00",X"A2",X"28",X"20",
		X"1D",X"D8",X"A9",X"00",X"A0",X"84",X"20",X"EF",X"D7",X"A9",X"00",X"20",X"10",X"D8",X"A0",X"00",
		X"AD",X"70",X"56",X"91",X"11",X"C8",X"AD",X"71",X"56",X"91",X"11",X"E6",X"11",X"E6",X"11",X"A9",
		X"01",X"20",X"10",X"D8",X"AD",X"C8",X"04",X"F0",X"0E",X"A2",X"02",X"20",X"B7",X"DC",X"AD",X"C9",
		X"04",X"18",X"69",X"01",X"20",X"AF",X"D7",X"A2",X"18",X"20",X"B7",X"DC",X"AD",X"22",X"04",X"20",
		X"A1",X"DC",X"48",X"4A",X"4A",X"4A",X"4A",X"38",X"20",X"AF",X"D7",X"68",X"29",X"0F",X"18",X"20",
		X"AF",X"D7",X"A2",X"12",X"20",X"B7",X"DC",X"A2",X"14",X"20",X"B7",X"DC",X"A2",X"1C",X"20",X"B7",
		X"DC",X"A9",X"90",X"A2",X"02",X"20",X"64",X"DC",X"A2",X"1E",X"20",X"B7",X"DC",X"A9",X"03",X"85",
		X"1E",X"AD",X"5D",X"04",X"38",X"E9",X"04",X"85",X"1D",X"A9",X"C8",X"85",X"1C",X"A5",X"1D",X"10",
		X"03",X"4C",X"38",X"DC",X"20",X"F9",X"D7",X"A9",X"BB",X"A6",X"1C",X"20",X"1D",X"D8",X"A0",X"C1",
		X"A5",X"1E",X"C9",X"02",X"D0",X"0D",X"A5",X"6F",X"4A",X"4A",X"29",X"07",X"D0",X"02",X"A9",X"07",
		X"09",X"E0",X"A8",X"A9",X"00",X"20",X"EF",X"D7",X"A5",X"1D",X"18",X"69",X"01",X"20",X"A1",X"DC",
		X"48",X"4A",X"4A",X"4A",X"4A",X"38",X"20",X"AF",X"D7",X"68",X"29",X"0F",X"18",X"20",X"AF",X"D7",
		X"A9",X"00",X"8D",X"37",X"04",X"8D",X"38",X"04",X"8D",X"39",X"04",X"A9",X"10",X"A2",X"00",X"20",
		X"1D",X"D8",X"A5",X"1D",X"F0",X"1D",X"4A",X"4A",X"38",X"E9",X"01",X"85",X"1B",X"0A",X"65",X"1B",
		X"AA",X"BD",X"24",X"DE",X"8D",X"37",X"04",X"BD",X"25",X"DE",X"8D",X"38",X"04",X"BD",X"26",X"DE",
		X"8D",X"39",X"04",X"AD",X"5D",X"04",X"C5",X"1D",X"D0",X"0C",X"AD",X"39",X"04",X"48",X"AD",X"38",
		X"04",X"48",X"AD",X"37",X"04",X"48",X"AD",X"37",X"04",X"4A",X"4A",X"4A",X"4A",X"38",X"F0",X"01",
		X"18",X"20",X"AF",X"D7",X"AD",X"37",X"04",X"20",X"60",X"DA",X"AD",X"38",X"04",X"4A",X"4A",X"4A",
		X"4A",X"20",X"60",X"DA",X"AD",X"38",X"04",X"29",X"0F",X"20",X"60",X"DA",X"AD",X"39",X"04",X"4A",
		X"4A",X"4A",X"4A",X"18",X"20",X"AF",X"D7",X"AD",X"39",X"04",X"18",X"20",X"AF",X"D7",X"20",X"F9",
		X"D7",X"A9",X"0C",X"A6",X"1C",X"20",X"1D",X"D8",X"A5",X"1D",X"29",X"78",X"4A",X"4A",X"C9",X"18",
		X"90",X"02",X"A9",X"16",X"AA",X"BD",X"58",X"DD",X"85",X"4C",X"BD",X"59",X"DD",X"85",X"4D",X"A9",
		X"FF",X"85",X"1B",X"E6",X"1B",X"A4",X"1B",X"B1",X"4C",X"A0",X"00",X"48",X"29",X"7F",X"AA",X"BD",
		X"C4",X"5D",X"91",X"11",X"C8",X"BD",X"C5",X"5D",X"91",X"11",X"A5",X"11",X"18",X"69",X"02",X"85",
		X"11",X"90",X"02",X"E6",X"12",X"68",X"10",X"DB",X"A5",X"1D",X"30",X"05",X"CD",X"2B",X"06",X"B0",
		X"13",X"18",X"69",X"04",X"85",X"1D",X"A5",X"1C",X"38",X"E9",X"0C",X"85",X"1C",X"C6",X"1E",X"F0",
		X"03",X"4C",X"2D",X"DB",X"68",X"8D",X"37",X"04",X"68",X"8D",X"38",X"04",X"68",X"8D",X"39",X"04",
		X"20",X"A2",X"D7",X"60",X"20",X"1D",X"D8",X"A0",X"C2",X"A9",X"00",X"20",X"EF",X"D7",X"A9",X"01",
		X"A8",X"20",X"10",X"D8",X"A9",X"16",X"AA",X"A9",X"2F",X"20",X"E3",X"D7",X"A0",X"87",X"A9",X"00",
		X"20",X"EF",X"D7",X"A9",X"00",X"AA",X"A9",X"2C",X"20",X"E3",X"D7",X"A0",X"00",X"A9",X"00",X"20",
		X"EF",X"D7",X"A9",X"01",X"20",X"10",X"D8",X"A9",X"10",X"A2",X"FE",X"A0",X"00",X"20",X"1D",X"D8",
		X"60",X"F8",X"85",X"19",X"A9",X"00",X"85",X"1B",X"A0",X"07",X"06",X"19",X"A5",X"1B",X"65",X"1B",
		X"85",X"1B",X"88",X"10",X"F5",X"D8",X"60",X"BD",X"29",X"E0",X"8E",X"02",X"03",X"85",X"1C",X"AC",
		X"02",X"03",X"B1",X"9B",X"85",X"9D",X"C8",X"B1",X"9B",X"85",X"9E",X"A0",X"00",X"B1",X"9D",X"85",
		X"1B",X"20",X"F9",X"D7",X"A9",X"00",X"85",X"0C",X"A9",X"01",X"20",X"10",X"D8",X"A5",X"1B",X"A6",
		X"1C",X"20",X"1D",X"D8",X"AC",X"02",X"03",X"B1",X"9B",X"85",X"9D",X"C8",X"B1",X"9B",X"85",X"9E",
		X"AE",X"02",X"03",X"BD",X"28",X"E0",X"48",X"4A",X"4A",X"4A",X"4A",X"09",X"C0",X"A8",X"29",X"08",
		X"F0",X"09",X"AD",X"D0",X"03",X"29",X"C0",X"D0",X"02",X"A0",X"00",X"A9",X"00",X"20",X"EF",X"D7",
		X"68",X"A0",X"10",X"29",X"0F",X"C9",X"01",X"F0",X"04",X"A0",X"68",X"A9",X"01",X"20",X"12",X"D8",
		X"A0",X"01",X"A9",X"00",X"85",X"1B",X"B1",X"9D",X"85",X"1C",X"29",X"7F",X"C8",X"84",X"1D",X"AA",
		X"BD",X"C4",X"5D",X"A4",X"1B",X"91",X"11",X"C8",X"BD",X"C5",X"5D",X"91",X"11",X"C8",X"84",X"1B",
		X"A4",X"1D",X"24",X"1C",X"10",X"E0",X"A4",X"1B",X"88",X"4C",X"05",X"D8",X"8E",X"02",X"03",X"85",
		X"1B",X"A9",X"00",X"85",X"1C",X"4C",X"D4",X"DC",X"70",X"DD",X"7F",X"DD",X"8E",X"DD",X"9D",X"DD",
		X"AC",X"DD",X"BB",X"DD",X"CA",X"DD",X"D9",X"DD",X"E8",X"DD",X"F7",X"DD",X"06",X"DE",X"15",X"DE",
		X"00",X"00",X"00",X"20",X"1E",X"38",X"00",X"3A",X"3E",X"38",X"1E",X"00",X"00",X"00",X"80",X"00",
		X"00",X"00",X"20",X"16",X"38",X"00",X"32",X"3E",X"3C",X"00",X"00",X"00",X"00",X"80",X"00",X"00",
		X"00",X"26",X"30",X"3C",X"1E",X"30",X"3A",X"1E",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",
		X"00",X"3E",X"30",X"38",X"1E",X"16",X"2C",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"16",
		X"42",X"1E",X"3A",X"32",X"2E",X"1E",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"26",
		X"30",X"3A",X"16",X"30",X"1E",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"3C",X"3E",X"18",
		X"3E",X"2C",X"16",X"38",X"00",X"00",X"00",X"00",X"80",X"3C",X"32",X"3C",X"16",X"2C",X"2C",X"46",
		X"00",X"16",X"42",X"1E",X"3A",X"32",X"2E",X"9E",X"2C",X"3E",X"30",X"16",X"3C",X"26",X"1A",X"00",
		X"20",X"38",X"26",X"30",X"22",X"1E",X"80",X"00",X"00",X"3C",X"32",X"00",X"3C",X"24",X"1E",X"00",
		X"2E",X"16",X"44",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"1A",X"32",X"3A",X"2E",X"26",X"1A",
		X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"30",X"32",X"00",X"42",X"16",X"46",X"00",
		X"00",X"00",X"00",X"80",X"02",X"50",X"00",X"05",X"00",X"00",X"07",X"50",X"00",X"10",X"00",X"00",
		X"12",X"50",X"00",X"15",X"00",X"00",X"17",X"50",X"00",X"21",X"50",X"00",X"25",X"50",X"00",X"29",
		X"50",X"00",X"33",X"50",X"00",X"37",X"50",X"00",X"41",X"50",X"00",X"45",X"50",X"00",X"49",X"50",
		X"00",X"53",X"50",X"00",X"57",X"50",X"00",X"61",X"50",X"00",X"65",X"50",X"00",X"69",X"50",X"00",
		X"73",X"50",X"00",X"77",X"50",X"00",X"81",X"50",X"00",X"85",X"50",X"00",X"89",X"50",X"00",X"A2",
		X"2C",X"20",X"B7",X"DC",X"A5",X"8C",X"29",X"03",X"D0",X"04",X"A9",X"02",X"D0",X"02",X"A5",X"8D",
		X"20",X"A1",X"DC",X"48",X"4A",X"4A",X"4A",X"4A",X"38",X"20",X"AF",X"D7",X"68",X"29",X"0F",X"18",
		X"20",X"AF",X"D7",X"A5",X"8C",X"29",X"03",X"49",X"03",X"D0",X"0C",X"A5",X"95",X"F0",X"08",X"A9",
		X"52",X"AA",X"A9",X"5F",X"20",X"E3",X"D7",X"60",X"88",X"E0",X"BA",X"E0",X"BA",X"E0",X"DC",X"E0",
		X"FE",X"E0",X"16",X"E1",X"74",X"E1",X"E1",X"E1",X"4E",X"E2",X"7D",X"E2",X"B6",X"E2",X"F5",X"E2",
		X"FB",X"E2",X"16",X"E3",X"31",X"E3",X"62",X"E3",X"93",X"E3",X"D4",X"E3",X"DE",X"E3",X"22",X"E4",
		X"63",X"E4",X"A8",X"E4",X"BA",X"E4",X"D6",X"E4",X"17",X"E5",X"51",X"E5",X"69",X"E5",X"8B",X"E5",
		X"D7",X"E5",X"B1",X"E5",X"00",X"E6",X"0E",X"E6",X"13",X"E6",X"1A",X"E6",X"1F",X"E6",X"2C",X"E6",
		X"49",X"E6",X"52",X"E6",X"62",X"E6",X"71",X"E6",X"8B",X"E6",X"A3",X"E6",X"B0",X"E6",X"BC",X"E6",
		X"C9",X"E6",X"E3",X"E6",X"02",X"E7",X"26",X"E7",X"92",X"E0",X"C2",X"E0",X"C2",X"E0",X"E8",X"E0",
		X"03",X"E1",X"2A",X"E1",X"8B",X"E1",X"FB",X"E1",X"67",X"E2",X"A0",X"E2",X"DF",X"E2",X"F5",X"E2",
		X"01",X"E3",X"1C",X"E3",X"4C",X"E3",X"7D",X"E3",X"A0",X"E3",X"D4",X"E3",X"ED",X"E3",X"30",X"E4",
		X"72",X"E4",X"A8",X"E4",X"BA",X"E4",X"E7",X"E4",X"2B",X"E5",X"57",X"E5",X"75",X"E5",X"9B",X"E5",
		X"EA",X"E5",X"C1",X"E5",X"00",X"E6",X"0E",X"E6",X"13",X"E6",X"1A",X"E6",X"1F",X"E6",X"2C",X"E6",
		X"49",X"E6",X"52",X"E6",X"62",X"E6",X"71",X"E6",X"8B",X"E6",X"A3",X"E6",X"B0",X"E6",X"BC",X"E6",
		X"C9",X"E6",X"E3",X"E6",X"02",X"E7",X"26",X"E7",X"A0",X"E0",X"CA",X"E0",X"CA",X"E0",X"EF",X"E0",
		X"09",X"E1",X"43",X"E1",X"AA",X"E1",X"16",X"E2",X"6E",X"E2",X"A7",X"E2",X"E6",X"E2",X"F5",X"E2",
		X"08",X"E3",X"24",X"E3",X"5B",X"E3",X"8C",X"E3",X"B6",X"E3",X"D4",X"E3",X"FF",X"E3",X"41",X"E4",
		X"84",X"E4",X"A8",X"E4",X"C3",X"E4",X"F6",X"E4",X"39",X"E5",X"5E",X"E5",X"7C",X"E5",X"A2",X"E5",
		X"F1",X"E5",X"C8",X"E5",X"00",X"E6",X"0E",X"E6",X"13",X"E6",X"1A",X"E6",X"1F",X"E6",X"2C",X"E6",
		X"49",X"E6",X"52",X"E6",X"62",X"E6",X"71",X"E6",X"8B",X"E6",X"A3",X"E6",X"B0",X"E6",X"BC",X"E6",
		X"C9",X"E6",X"E3",X"E6",X"02",X"E7",X"26",X"E7",X"AA",X"E0",X"D3",X"E0",X"D3",X"E0",X"F6",X"E0",
		X"0F",X"E1",X"60",X"E1",X"C4",X"E1",X"31",X"E2",X"75",X"E2",X"AE",X"E2",X"ED",X"E2",X"F5",X"E2",
		X"0E",X"E3",X"2A",X"E3",X"53",X"E3",X"84",X"E3",X"C5",X"E3",X"D4",X"E3",X"10",X"E4",X"52",X"E4",
		X"96",X"E4",X"A8",X"E4",X"CC",X"E4",X"07",X"E5",X"45",X"E5",X"63",X"E5",X"83",X"E5",X"A9",X"E5");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
