library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_VEC_ROM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_VEC_ROM_1 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"B9",X"00",X"02",X"29",X"3C",X"4A",X"4A",X"AA",X"BD",X"F8",X"02",X"10",X"31",X"86",X"1A",X"A9",
		X"05",X"20",X"B2",X"48",X"20",X"50",X"6D",X"EE",X"E7",X"02",X"B9",X"00",X"02",X"48",X"20",X"EB",
		X"61",X"68",X"9D",X"00",X"02",X"A9",X"00",X"99",X"00",X"02",X"A6",X"1A",X"BD",X"F8",X"02",X"10",
		X"1D",X"48",X"A9",X"7F",X"9D",X"F8",X"02",X"68",X"4A",X"29",X"0F",X"AA",X"10",X"EE",X"4A",X"B0",
		X"10",X"A9",X"00",X"9D",X"F8",X"02",X"A9",X"20",X"20",X"B2",X"48",X"20",X"AC",X"49",X"A6",X"0E",
		X"60",X"A9",X"10",X"86",X"1A",X"20",X"B2",X"48",X"20",X"50",X"6D",X"20",X"EB",X"61",X"EE",X"E7",
		X"02",X"EE",X"FF",X"02",X"A5",X"1A",X"0A",X"0A",X"09",X"42",X"9D",X"00",X"02",X"86",X"10",X"A6",
		X"1A",X"A9",X"7E",X"9D",X"F8",X"02",X"A5",X"79",X"69",X"20",X"9D",X"F1",X"02",X"20",X"A7",X"48",
		X"86",X"1A",X"A6",X"10",X"20",X"52",X"6D",X"20",X"EB",X"61",X"EE",X"E7",X"02",X"A5",X"1A",X"0A",
		X"0A",X"09",X"42",X"9D",X"00",X"02",X"A6",X"1A",X"A9",X"7E",X"9D",X"F8",X"02",X"A5",X"79",X"E9",
		X"20",X"9D",X"F1",X"02",X"A6",X"0E",X"60",X"A2",X"06",X"BD",X"F8",X"02",X"F0",X"03",X"CA",X"10",
		X"F8",X"60",X"A6",X"0E",X"F0",X"04",X"E0",X"04",X"90",X"F7",X"18",X"4C",X"44",X"6C",X"86",X"10",
		X"A0",X"19",X"84",X"11",X"E6",X"19",X"BD",X"00",X"02",X"4A",X"4A",X"29",X"0F",X"AA",X"BC",X"F8",
		X"02",X"C0",X"04",X"90",X"1C",X"A5",X"76",X"29",X"0F",X"D0",X"07",X"98",X"38",X"E9",X"02",X"9D",
		X"F8",X"02",X"AD",X"19",X"02",X"F0",X"02",X"10",X"0A",X"98",X"29",X"01",X"09",X"02",X"9D",X"F8",
		X"02",X"E6",X"11",X"A4",X"11",X"86",X"1A",X"A6",X"10",X"20",X"22",X"4A",X"20",X"FD",X"49",X"85",
		X"13",X"A5",X"0C",X"85",X"12",X"A5",X"11",X"18",X"69",X"21",X"A8",X"8A",X"69",X"21",X"AA",X"20",
		X"22",X"4A",X"20",X"FD",X"49",X"20",X"32",X"4A",X"A6",X"1A",X"85",X"12",X"A0",X"19",X"C4",X"11",
		X"D0",X"19",X"49",X"80",X"E5",X"79",X"10",X"02",X"49",X"FF",X"C9",X"10",X"B0",X"0D",X"A5",X"12",
		X"FD",X"F1",X"02",X"10",X"02",X"49",X"FF",X"C9",X"40",X"90",X"31",X"A5",X"12",X"38",X"FD",X"F1",
		X"02",X"85",X"12",X"10",X"02",X"49",X"FF",X"C9",X"08",X"90",X"21",X"A9",X"01",X"A0",X"19",X"C4",
		X"11",X"D0",X"0D",X"A6",X"19",X"E0",X"07",X"90",X"02",X"A2",X"00",X"BD",X"A4",X"49",X"A6",X"1A",
		X"06",X"12",X"90",X"02",X"49",X"FF",X"7D",X"F1",X"02",X"9D",X"F1",X"02",X"AD",X"F0",X"02",X"4A",
		X"18",X"65",X"D3",X"0A",X"CD",X"57",X"69",X"90",X"03",X"AD",X"57",X"69",X"6D",X"58",X"69",X"85",
		X"11",X"48",X"BD",X"F1",X"02",X"20",X"FE",X"70",X"20",X"BB",X"49",X"A6",X"10",X"9D",X"21",X"02",
		X"68",X"85",X"11",X"A6",X"1A",X"BD",X"F1",X"02",X"20",X"01",X"71",X"20",X"BB",X"49",X"A6",X"10",
		X"9D",X"42",X"02",X"60",X"01",X"02",X"03",X"03",X"03",X"04",X"04",X"11",X"CE",X"FF",X"02",X"D0",
		X"09",X"98",X"48",X"A0",X"3F",X"20",X"16",X"77",X"68",X"A8",X"60",X"A8",X"10",X"05",X"49",X"FF",
		X"18",X"69",X"01",X"85",X"12",X"A9",X"00",X"85",X"13",X"06",X"11",X"B0",X"0D",X"D0",X"12",X"A5",
		X"13",X"C0",X"00",X"10",X"04",X"49",X"FF",X"69",X"00",X"60",X"A5",X"13",X"18",X"65",X"12",X"85",
		X"13",X"46",X"12",X"D0",X"E4",X"F0",X"E8",X"C9",X"10",X"90",X"11",X"C9",X"F0",X"B0",X"0D",X"85",
		X"15",X"A9",X"00",X"38",X"E5",X"0C",X"85",X"0C",X"A9",X"00",X"E5",X"15",X"60",X"C9",X"04",X"90",
		X"FB",X"C9",X"FC",X"B0",X"F7",X"A4",X"D3",X"C0",X"05",X"90",X"DC",X"A4",X"19",X"C0",X"03",X"90",
		X"D6",X"85",X"15",X"8A",X"E0",X"21",X"B0",X"01",X"4A",X"4A",X"6A",X"45",X"15",X"30",X"D2",X"A5",
		X"15",X"60",X"B9",X"A5",X"02",X"38",X"FD",X"A5",X"02",X"85",X"0C",X"B9",X"63",X"02",X"FD",X"63",
		X"02",X"60",X"85",X"14",X"10",X"03",X"20",X"B6",X"70",X"85",X"15",X"A5",X"13",X"10",X"03",X"20",
		X"B6",X"70",X"05",X"15",X"A2",X"07",X"0A",X"30",X"03",X"CA",X"D0",X"FA",X"E0",X"04",X"B0",X"12",
		X"46",X"13",X"66",X"12",X"46",X"14",X"66",X"0C",X"CA",X"10",X"F5",X"A6",X"12",X"A4",X"0C",X"4C",
		X"9E",X"70",X"06",X"12",X"26",X"13",X"06",X"0C",X"26",X"14",X"E8",X"E0",X"07",X"90",X"F3",X"A6",
		X"13",X"A4",X"14",X"B0",X"EA",X"4A",X"4A",X"4A",X"29",X"0F",X"AA",X"BD",X"F8",X"02",X"4A",X"A9",
		X"00",X"6A",X"6A",X"85",X"11",X"BD",X"F1",X"02",X"4A",X"4A",X"24",X"11",X"50",X"02",X"29",X"1E",
		X"29",X"3E",X"05",X"11",X"A8",X"BE",X"2B",X"50",X"B9",X"2A",X"50",X"4C",X"D5",X"7C",X"AD",X"F0",
		X"02",X"F0",X"13",X"18",X"A2",X"02",X"69",X"02",X"C9",X"05",X"90",X"03",X"E8",X"A9",X"05",X"86",
		X"11",X"CD",X"E7",X"02",X"B0",X"01",X"60",X"AE",X"FF",X"02",X"D0",X"FA",X"AC",X"E7",X"02",X"BD",
		X"00",X"02",X"D0",X"02",X"86",X"10",X"10",X"01",X"88",X"E8",X"E0",X"19",X"90",X"F1",X"A6",X"1E",
		X"B5",X"D1",X"F0",X"04",X"C4",X"11",X"90",X"DE",X"A0",X"1A",X"94",X"D1",X"A6",X"10",X"20",X"E7",
		X"69",X"20",X"4D",X"4B",X"A0",X"02",X"84",X"DD",X"98",X"0A",X"0A",X"09",X"42",X"9D",X"00",X"02",
		X"EE",X"E7",X"02",X"EE",X"FF",X"02",X"B9",X"47",X"4B",X"99",X"F8",X"02",X"B9",X"4A",X"4B",X"99",
		X"F1",X"02",X"B9",X"3B",X"4B",X"18",X"7D",X"A5",X"02",X"9D",X"A5",X"02",X"B9",X"3E",X"4B",X"7D",
		X"63",X"02",X"9D",X"63",X"02",X"B9",X"41",X"4B",X"18",X"7D",X"C6",X"02",X"9D",X"C6",X"02",X"B9",
		X"44",X"4B",X"7D",X"84",X"02",X"9D",X"84",X"02",X"88",X"30",X"8B",X"86",X"10",X"20",X"52",X"6D",
		X"84",X"11",X"A4",X"10",X"20",X"EB",X"61",X"A4",X"11",X"10",X"AD",X"00",X"58",X"70",X"00",X"FF",
		X"00",X"40",X"50",X"00",X"FF",X"00",X"00",X"83",X"85",X"81",X"F0",X"98",X"40",X"20",X"53",X"4B",
		X"9D",X"21",X"02",X"A0",X"06",X"AD",X"0A",X"2C",X"10",X"02",X"A0",X"FA",X"98",X"9D",X"42",X"02",
		X"60",X"00",X"03",X"06",X"09",X"0C",X"10",X"13",X"16",X"19",X"1C",X"1F",X"22",X"25",X"28",X"2B",
		X"2E",X"31",X"33",X"36",X"39",X"3C",X"3F",X"41",X"44",X"47",X"49",X"4C",X"4E",X"51",X"53",X"55",
		X"58",X"5A",X"5C",X"5E",X"60",X"62",X"64",X"66",X"68",X"6A",X"6B",X"6D",X"6F",X"70",X"71",X"73",
		X"74",X"75",X"76",X"78",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"7F",X"7F",X"A5",X"76",X"29",X"03",X"AA",X"18",X"69",X"FE",X"75",X"86",X"95",X"86",X"29",X"F0",
		X"18",X"75",X"86",X"0A",X"20",X"C6",X"6E",X"B9",X"02",X"50",X"85",X"10",X"B9",X"03",X"50",X"85",
		X"11",X"8A",X"0A",X"AA",X"0A",X"29",X"04",X"45",X"09",X"85",X"09",X"BD",X"9D",X"77",X"0A",X"85",
		X"03",X"BD",X"9E",X"77",X"2A",X"49",X"C0",X"85",X"04",X"A2",X"0C",X"20",X"21",X"62",X"4C",X"D6",
		X"79",X"A5",X"22",X"F0",X"0E",X"A5",X"74",X"D0",X"03",X"4C",X"F6",X"4C",X"C6",X"74",X"20",X"EB",
		X"60",X"18",X"60",X"85",X"13",X"A5",X"8D",X"29",X"03",X"D0",X"06",X"A9",X"02",X"85",X"8C",X"D0",
		X"56",X"18",X"69",X"07",X"A8",X"A5",X"42",X"25",X"43",X"10",X"4C",X"20",X"59",X"71",X"A5",X"8C",
		X"C9",X"40",X"B0",X"FE",X"85",X"10",X"A0",X"0B",X"20",X"59",X"71",X"A2",X"00",X"86",X"11",X"E8",
		X"86",X"12",X"F8",X"46",X"10",X"90",X"07",X"A5",X"11",X"18",X"65",X"12",X"85",X"11",X"F0",X"08",
		X"A5",X"12",X"65",X"12",X"85",X"12",X"90",X"EB",X"D8",X"A2",X"00",X"A0",X"01",X"A9",X"11",X"38",
		X"20",X"95",X"7C",X"A5",X"8D",X"29",X"03",X"C9",X"03",X"D0",X"0C",X"A5",X"8F",X"4A",X"90",X"07",
		X"A9",X"20",X"A2",X"CB",X"20",X"D5",X"7C",X"A0",X"06",X"A6",X"8C",X"D0",X"02",X"86",X"8A",X"AD",
		X"01",X"28",X"4A",X"90",X"10",X"24",X"8A",X"30",X"0C",X"E0",X"01",X"90",X"04",X"D0",X"06",X"66",
		X"13",X"A0",X"0C",X"D0",X"08",X"A9",X"FF",X"85",X"8A",X"C0",X"0C",X"D0",X"09",X"20",X"DB",X"60",
		X"18",X"A9",X"00",X"85",X"85",X"60",X"8A",X"F0",X"F7",X"20",X"DB",X"60",X"A4",X"8C",X"A2",X"01",
		X"AD",X"03",X"24",X"30",X"20",X"C0",X"02",X"90",X"49",X"AD",X"04",X"24",X"10",X"44",X"8D",X"04",
		X"3C",X"20",X"D0",X"60",X"20",X"E3",X"7B",X"20",X"59",X"69",X"20",X"1B",X"6A",X"A5",X"6E",X"85",
		X"70",X"A2",X"02",X"C6",X"8C",X"86",X"22",X"C6",X"8C",X"8E",X"04",X"3C",X"86",X"85",X"20",X"D0",
		X"60",X"20",X"E3",X"7B",X"20",X"1B",X"6A",X"A9",X"80",X"85",X"74",X"0A",X"85",X"1E",X"85",X"1F",
		X"85",X"20",X"85",X"9A",X"85",X"99",X"A5",X"6E",X"85",X"6F",X"A9",X"04",X"85",X"84",X"8D",X"00",
		X"3E",X"60",X"A5",X"76",X"29",X"0F",X"D0",X"0C",X"A9",X"01",X"C5",X"8C",X"F0",X"02",X"A9",X"03",
		X"45",X"85",X"85",X"85",X"18",X"60",X"A5",X"76",X"29",X"3F",X"D0",X"0A",X"AD",X"ED",X"02",X"C9",
		X"08",X"F0",X"03",X"CE",X"ED",X"02",X"A6",X"1E",X"B5",X"6F",X"D0",X"1C",X"AD",X"1D",X"02",X"0D",
		X"1E",X"02",X"0D",X"1F",X"02",X"0D",X"20",X"02",X"D0",X"0E",X"A0",X"07",X"20",X"59",X"71",X"A5",
		X"22",X"C9",X"02",X"90",X"03",X"20",X"EB",X"60",X"AD",X"19",X"02",X"D0",X"37",X"AD",X"EB",X"02",
		X"C9",X"80",X"D0",X"30",X"A9",X"10",X"20",X"00",X"63",X"A6",X"22",X"A5",X"6F",X"05",X"70",X"F0",
		X"25",X"20",X"EB",X"67",X"CA",X"F0",X"1D",X"A9",X"80",X"85",X"74",X"A5",X"1E",X"49",X"01",X"AA",
		X"B5",X"6F",X"F0",X"10",X"86",X"1E",X"8A",X"6A",X"6A",X"8D",X"04",X"3C",X"8A",X"0A",X"85",X"1F",
		X"05",X"1E",X"85",X"20",X"18",X"60",X"86",X"21",X"A9",X"FF",X"85",X"22",X"A9",X"03",X"85",X"85",
		X"8D",X"04",X"3C",X"D0",X"EF",X"10",X"05",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"15",X"C7",X"FA",X"C6",X"DB",X"C6",X"C4",X"C6",X"0D",X"F8",X"78",X"F8",X"0D",X"FD",X"78",X"F8",
		X"09",X"FD",X"78",X"F8",X"0B",X"F1",X"78",X"F8",X"0A",X"F5",X"78",X"F8",X"08",X"F9",X"78",X"F8",
		X"09",X"F3",X"78",X"F8",X"0D",X"F3",X"78",X"F8",X"80",X"54",X"00",X"06",X"78",X"F8",X"0F",X"F1",
		X"78",X"F8",X"0A",X"FE",X"00",X"D0",X"00",X"30",X"80",X"07",X"78",X"F8",X"80",X"37",X"80",X"07",
		X"78",X"F8",X"80",X"37",X"80",X"03",X"78",X"F8",X"E0",X"40",X"A0",X"02",X"78",X"F8",X"C0",X"35",
		X"80",X"03",X"78",X"F8",X"80",X"33",X"00",X"00",X"78",X"F8",X"A0",X"42",X"E0",X"00",X"78",X"F8",
		X"A0",X"42",X"E0",X"04",X"78",X"F8",X"E0",X"44",X"80",X"07",X"78",X"F8",X"E0",X"40",X"A0",X"06",
		X"78",X"F8",X"00",X"D0",X"07",X"F8",X"78",X"F8",X"07",X"FF",X"78",X"F8",X"03",X"FF",X"78",X"F8",
		X"C0",X"40",X"40",X"02",X"78",X"F8",X"80",X"35",X"00",X"03",X"78",X"F8",X"00",X"FB",X"78",X"F8",
		X"40",X"42",X"C0",X"00",X"78",X"F8",X"40",X"42",X"C0",X"04",X"78",X"F8",X"C0",X"44",X"00",X"07",
		X"78",X"F8",X"C0",X"40",X"40",X"06",X"78",X"F8",X"00",X"D0",X"00",X"30",X"80",X"06",X"78",X"F8",
		X"80",X"36",X"80",X"06",X"78",X"F8",X"80",X"36",X"80",X"02",X"78",X"F8",X"40",X"31",X"C0",X"03",
		X"78",X"F8",X"40",X"35",X"80",X"02",X"78",X"F8",X"80",X"32",X"00",X"00",X"78",X"F8",X"C0",X"33",
		X"40",X"01",X"78",X"F8",X"C0",X"33",X"40",X"05",X"78",X"F8",X"A0",X"44",X"80",X"06",X"78",X"F8",
		X"40",X"31",X"C0",X"07",X"78",X"F8",X"00",X"D0",X"0E",X"F1",X"CA",X"F8",X"0B",X"F6",X"00",X"60",
		X"80",X"D6",X"DB",X"F6",X"CA",X"F8",X"DB",X"F2",X"DF",X"F2",X"CD",X"F2",X"CD",X"F8",X"CD",X"F6",
		X"DF",X"F6",X"00",X"D0",X"09",X"F0",X"7B",X"F1",X"78",X"F1",X"7F",X"F2",X"7F",X"F0",X"79",X"F6",
		X"7E",X"F8",X"78",X"F7",X"7B",X"F7",X"7B",X"F1",X"79",X"F5",X"79",X"F9",X"7F",X"F2",X"80",X"30",
		X"00",X"02",X"80",X"41",X"C0",X"72",X"00",X"32",X"80",X"74",X"60",X"41",X"40",X"77",X"A0",X"44",
		X"00",X"77",X"80",X"37",X"C0",X"72",X"C0",X"44",X"E0",X"77",X"00",X"47",X"80",X"70",X"60",X"46",
		X"A0",X"73",X"A0",X"41",X"C0",X"72",X"80",X"35",X"40",X"72",X"60",X"42",X"A0",X"71",X"60",X"41",
		X"60",X"77",X"80",X"21",X"80",X"03",X"20",X"42",X"80",X"72",X"80",X"23",X"00",X"76",X"C0",X"40",
		X"80",X"77",X"40",X"45",X"C0",X"76",X"C0",X"36",X"40",X"73",X"A0",X"45",X"A0",X"77",X"C0",X"46",
		X"20",X"71",X"A0",X"45",X"E0",X"73",X"20",X"42",X"80",X"72",X"00",X"35",X"80",X"72",X"80",X"42",
		X"20",X"71",X"C0",X"40",X"A0",X"77",X"00",X"22",X"80",X"03",X"80",X"42",X"E0",X"71",X"80",X"23",
		X"00",X"76",X"00",X"40",X"A0",X"77",X"A0",X"45",X"80",X"76",X"40",X"36",X"C0",X"73",X"40",X"46",
		X"40",X"77",X"80",X"46",X"A0",X"71",X"60",X"54",X"10",X"72",X"60",X"42",X"00",X"72",X"80",X"34",
		X"C0",X"72",X"C0",X"42",X"80",X"70",X"00",X"40",X"80",X"77",X"03",X"F3",X"C0",X"42",X"60",X"71",
		X"77",X"F3",X"C0",X"44",X"80",X"77",X"20",X"46",X"20",X"76",X"A0",X"44",X"20",X"72",X"E0",X"46",
		X"E0",X"76",X"20",X"46",X"20",X"72",X"00",X"50",X"20",X"72",X"E0",X"42",X"80",X"71",X"00",X"30",
		X"C0",X"72",X"C0",X"42",X"00",X"70",X"A0",X"44",X"80",X"77",X"80",X"23",X"00",X"02",X"00",X"43",
		X"E0",X"70",X"00",X"22",X"80",X"77",X"60",X"45",X"40",X"77",X"80",X"46",X"A0",X"75",X"40",X"44",
		X"20",X"72",X"40",X"47",X"40",X"76",X"C0",X"45",X"80",X"72",X"70",X"50",X"20",X"72",X"00",X"43",
		X"C0",X"70",X"C0",X"30",X"C0",X"72",X"C0",X"42",X"80",X"74",X"60",X"45",X"60",X"77",X"80",X"23",
		X"80",X"01",X"40",X"43",X"40",X"70",X"C0",X"30",X"00",X"76",X"7F",X"F6",X"E0",X"46",X"20",X"75",
		X"40",X"40",X"40",X"72",X"C0",X"47",X"80",X"75",X"20",X"45",X"C0",X"72",X"A0",X"41",X"E0",X"73",
		X"20",X"43",X"40",X"70",X"40",X"31",X"C0",X"72",X"80",X"42",X"20",X"75",X"7F",X"F6",X"00",X"32",
		X"80",X"00",X"20",X"43",X"80",X"74",X"00",X"21",X"80",X"77",X"A0",X"46",X"A0",X"76",X"E0",X"46",
		X"A0",X"74",X"80",X"40",X"40",X"72",X"E0",X"47",X"C0",X"74",X"A0",X"44",X"E0",X"72",X"60",X"42",
		X"80",X"73",X"20",X"43",X"60",X"74",X"80",X"31",X"80",X"72",X"60",X"42",X"A0",X"75",X"80",X"46");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
