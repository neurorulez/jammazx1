-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "9797979349294A02942528493FE22AAA6AAAAA712E050080A16135DFDEA3B3FD";
    attribute INIT_01 of inst : label is "210130DF1E20023FBA010DB67915D4929A4CC000CE6575AA0AA098CE19679797";
    attribute INIT_02 of inst : label is "B4E1150552009416A045530284C0AA502861184C1B6A126C39272882019A4C9B";
    attribute INIT_03 of inst : label is "F336492C92A3A8EDD893242211518A8C7473A39127F6F4ADF0521F62B642CFA8";
    attribute INIT_04 of inst : label is "8454F77EE5B7DE7BFDF79EBF79E7BFDE79EBE12ED77000888888888888C44091";
    attribute INIT_05 of inst : label is "D7780F5FBFC804C965E135DA64D4449A9B06CB0F616C3FDE7D6DBB4959FE610A";
    attribute INIT_06 of inst : label is "000000088A288D162202DB9B9412B26B27D8093E3684542D88C102143D94A466";
    attribute INIT_07 of inst : label is "51555DD75D15754D35F17499A1F753B9DD4EE6753B9D365994F97F9C9EC09000";
    attribute INIT_08 of inst : label is "659EDC202C2305140892CD7111149213D6021414004400057695959594D30D35";
    attribute INIT_09 of inst : label is "224898811188A281205D204965B67D892006252311BC8A08A3499514502C565D";
    attribute INIT_0A of inst : label is "94964CF5830DB364F649332D880317301810AAAAAAAACB301000189DF5B34000";
    attribute INIT_0B of inst : label is "32CEB30C80AF6ED6AB76B4F59BF6B75FB5A7AEDBB5AADDAD3D66FDADD7ED69EB";
    attribute INIT_0C of inst : label is "A6B624B0A26D437EE1BBDA1088569484961049286FC62632202E41006800FAEA";
    attribute INIT_0D of inst : label is "DA86FF81B621BF96C377B42120B4A424B0E249437FE18D261B7D4F0DDC98C486";
    attribute INIT_0E of inst : label is "118A45809C2288D40031DE781E0781E000C6EEDF33A7B332B332802F5B125844";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000B6DB6DA4ECDC897";
    attribute INIT_10 of inst : label is "A4E8C49286FEA665BCEE8CA380CEEC63CC718BACBA87AE967F6B0924B9CA2E19";
    attribute INIT_11 of inst : label is "7B89B50DFDCCC7F4992D18D210DFD449286FEA665F36E8C4DA86FEE663A54D37";
    attribute INIT_12 of inst : label is "9373DC3814484F4677755552AA9D4E9D145D504A5454BA70A3DE6DDAD18DB61B";
    attribute INIT_13 of inst : label is "27FBB8C0B53249B376D9376D935BA534FB22EE4EEE11E04F8D0F8D0B890B890B";
    attribute INIT_14 of inst : label is "9F7E3EFC7DF8FBF1B7E36FC32A282FDF1FBE3F7C7EF8DDF1BBE40714572B88F6";
    attribute INIT_15 of inst : label is "000164220408102045D775873B2E31DD61CECB8C1B6C28A6AC312D60A44CD99B";
    attribute INIT_16 of inst : label is "8A00005E05A398CC662918C462316AB1CE64722294A3234414A55B6D24888800";
    attribute INIT_17 of inst : label is "6E2659DB899776E2659DB899758319491754D7473D673D773D673D7784417C11";
    attribute INIT_18 of inst : label is "D9303FBA418D6B041A028592A76432C10680A1A724975102A32635464C59A5FF";
    attribute INIT_19 of inst : label is "DD0F8713107B49524E3A66186227F18F989DFB1761BB9264A2945B640EE8A516";
    attribute INIT_1A of inst : label is "9624962494490D53BBBA22227274D34D34B61B9BB92486EDC60588282B5AD04D";
    attribute INIT_1B of inst : label is "A302C714D55464CAA8C9932AA3264EAA8C993AAA3264E3F363271DD3D8EBC824";
    attribute INIT_1C of inst : label is "0DDF7030B191316E0A0AAA32635464C58D5193161B9CB7186EE4921BB260632B";
    attribute INIT_1D of inst : label is "2DC61BB92486EE9819CEE8D0B5C535551932AA3264EAA8C9938FCC538C377B49";
    attribute INIT_1E of inst : label is "BC20444194F3E30DDED24377DC0C2C6444598282AA8C98D51931635464C586E7";
    attribute INIT_1F of inst : label is "C00000000000000000000000039009E339662013847AEE40278CE598804E11EB";
    attribute INIT_20 of inst : label is "90E91A0617742BC23287640ED650CE054AC21D68872FCC2AAA44F9FA7FCCF6C9";
    attribute INIT_21 of inst : label is "0AD3D1091E8DD34900103CB6A261427CA794EF24E04C2784BB498DD152E3A8E8";
    attribute INIT_22 of inst : label is "48971A4A829D6215A3744A0A0C42B468A8E89C38D68E886BA4DA3A258D146243";
    attribute INIT_23 of inst : label is "9921D11CA0645155FA1717F8045A114802381887C327420A8819410440230C4C";
    attribute INIT_24 of inst : label is "C22E91921061236B5293739E8903CCDAD4A49CE19207997EBE6DF72133327324";
    attribute INIT_25 of inst : label is "93C964B2391C8E4BA1D1E8F47A1861861854BBBBBB222222758B7DDD6FB3A36E";
    attribute INIT_26 of inst : label is "BC90B288E228B17A64AE1C6EA2C99649243D2C33164924924BB6D2486490E190";
    attribute INIT_27 of inst : label is "A0BD92C9AFE7DE4A64A1BDD2E9F3FA5FA509EC967CC95C940C9E4A8B0B772B2D";
    attribute INIT_28 of inst : label is "B25970774BA74BA15D92C992C85674BA74BA15D92C992C85674BBE066DFF4B74";
    attribute INIT_29 of inst : label is "B22C27D3B9E81FF6B8E7EDDFC070C63DBCF8D73E3FF5203CD7B9FCF1325935F7";
    attribute INIT_2A of inst : label is "CD34D864F2E0B48FBDB556D67EE11EF2BFC79DFF40C1A1081D3CCFB5624F9505";
    attribute INIT_2B of inst : label is "DA024279E7AAB4401F00C4A1F6D7FF7F032742EA7E01446294D80550004A5451";
    attribute INIT_2C of inst : label is "5CE811A67508D33A6CE24DBDD85C77425B3F3E6AFD3F865F7A68AE2E2B7C5638";
    attribute INIT_2D of inst : label is "A29A483050BDA8F6EE05B6B800007FFB62BA9CCDD33B0C98AAE74533AA99DA23";
    attribute INIT_2E of inst : label is "7F8FFBBF0A5D362F9ADD2E3BF686E359E648D6C7BF5971A7FCF5D33B0EA2A2A2";
    attribute INIT_2F of inst : label is "400000000000000002B33F5D4FD75375D4FD753EB53FFC850FA58576EEEEEEEB";
    attribute INIT_30 of inst : label is "0D31030008032003A6AE45191E25EF5596E1F897BD56E1D59F4251082B089A09";
    attribute INIT_31 of inst : label is "9215E0E8022044088150A3008C4208A8A71DD040404E007FCEE8200650214127";
    attribute INIT_32 of inst : label is "1DA91D00182051EA0190C1604CC00026535CEF964789DC600CA0C1158085921B";
    attribute INIT_33 of inst : label is "41F9FDFFD114662E62C444019F8BF1500C22E7A8001F188B89414787A2FAB333";
    attribute INIT_34 of inst : label is "00000101F4516E00000000020000000C0000009001000000001C550467F2AF15";
    attribute INIT_35 of inst : label is "33FFFFFF4927D3A76F400000000090080C30030E00007000024803C3EFF00000";
    attribute INIT_36 of inst : label is "DCF5D4000235F017FDF55DFDBD74FA4927FFFFFE633EE74E9FDF07F7DD3A7DC6";
    attribute INIT_37 of inst : label is "AE6540B4023E6A177028E9388E90A61F61D4F1F1C000F4E0F8C5C2ABDCD1393D";
    attribute INIT_38 of inst : label is "751D4741D0761D07C7FEC1FEB87FAA5FFF2EA97A41E9077D3B49DF6EDDBF705A";
    attribute INIT_39 of inst : label is "A7569DF6EFDB81CCCE4A77D3B53D1A9C06193D507672AAE4E551D9E029F2F9D4";
    attribute INIT_3A of inst : label is "A1958850FFF50078F001FEF17C3DDFBF800F00001E3FBFD50FFA87F6A5FBF2EF";
    attribute INIT_3B of inst : label is "4DCDE4264B944EB0BA0124C521442424000000000C000C004C4100000AA0A803";
    attribute INIT_3C of inst : label is "00000000122AA2D351A6A54D4772AA884128A21031C44411114A522294A44529";
    attribute INIT_3D of inst : label is "FFF1C01BFFEB8AA70F470D6E26AE349C5B1CD1B8D6BFD76337FAEC64B4023E6A";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000077D38027FFC7006FFFAE009";
    attribute INIT_3F of inst : label is "D000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "ADE5ADE0024FDF5FBE9F7D00802643334CCCCC29F2162C04B3289E7E7E66E3F7";
    attribute INIT_01 of inst : label is "63AD7C2502529340016CB26425B200240C999B6D99DA40145145111C8095ADE5";
    attribute INIT_02 of inst : label is "4E5FEB53A9CF9FBCDAFDA437D53BFF73FF6577A8043A6E5A8DC36DB0AABF5E23";
    attribute INIT_03 of inst : label is "0846C92592DCED326C2CD949E6223113888C449B3774EBD697F7B104473EBFEE";
    attribute INIT_04 of inst : label is "6EA49203392920AE165829C5960AF12482980B2480A000808080808080F93D9F";
    attribute INIT_05 of inst : label is "D2645BEADA82C92C9F4E4D24A9A99D3562F192D45E8B4349861926868464085D";
    attribute INIT_06 of inst : label is "C8C8C8C401040003497FE431BB7FB36B6C95A769EDBE9F6ED4C2F4CBE1D75ACE";
    attribute INIT_07 of inst : label is "EBBEF26D36DB4D3EFBCF0E314458A423A2900E9A423E44DE28333FA19F3CB288";
    attribute INIT_08 of inst : label is "DB289193CF8F25AFA8B24D2ACA414DF8F8000155112708B040228282802BEEBB";
    attribute INIT_09 of inst : label is "4981A75B415CB5F51449BB5925B2C955DB7D5ADC4132D3ED0253EDE6DA8BA906";
    attribute INIT_0A of inst : label is "DB99E55D75D0004AA4928CD979F6419DB5B27FFFFFFFBE767DBDB21D25964000";
    attribute INIT_0B of inst : label is "6C799641FF42BD4BF5CA4D596D5ACDEAD66AC9AB52ED5293564B76B3FBB59AB2";
    attribute INIT_0C of inst : label is "5949CB063593B090D84027396569293B21C29272020C8CA56D72D36A0EAE40B8";
    attribute INIT_0D of inst : label is "6F6120F2DBD84C7B3080DC62CA5B5BD90E34B79010DED2DC80C3B6402371892B";
    attribute INIT_0E of inst : label is "8339CDB3E308D11AEFA52F3D2F4BD2F4F62C9320B54846EECAC52A81ADE5830B";
    attribute INIT_0F of inst : label is "80000000000000000000000000000000000000000000000006DB6DB6DDBB004E";
    attribute INIT_10 of inst : label is "C997892520200A0C10B50B42509333302604C2C80CE84B24C886404126296983";
    attribute INIT_11 of inst : label is "C116DAC24094384B76D2D12DE4060896D20204A0A249B38B2561200A1A71B240";
    attribute INIT_12 of inst : label is "780532D22FC380AA0CFFFFFDFF92E1365A81DACA2FD9A4E46725B76D6516DD84";
    attribute INIT_13 of inst : label is "0A4ECC7F4F84B2EED9F66CBF2A0EEEC922C91114197F1B3A7878FAFA7878FAFA";
    attribute INIT_14 of inst : label is "51ADE1D946B787655ADE9D90F65F696AF274A5ABC9D2B6AF674EA12F8581624B";
    attribute INIT_15 of inst : label is "232393C448B322CD5A24D975E6C9AD324D3992E9565AC34CCB664A2DAFA9032E";
    attribute INIT_16 of inst : label is "3CC9C8B79E4CE330B8F2E31B84C795617E97D49B0BB5C5B9D85DE4B2F9131323";
    attribute INIT_17 of inst : label is "9188D2E4E274B9188D6E4E27582AD2E640D9A493D24BD64BD25BD6593726DE26";
    attribute INIT_18 of inst : label is "72D2A0459BDEF724D56D6927CE49F9CB355B5AD7386ABEF81CC8B03991761E3B";
    attribute INIT_19 of inst : label is "32934F8C3304FC109956A0D25A49082225C444B8C800248B2724E4C8A809C939";
    attribute INIT_1A of inst : label is "2D2B3D2B3E567EF84C4C4C4C04C96CB25B596480024B6111D1AE6D73F0F79F34";
    attribute INIT_1B of inst : label is "E8B72FB9B803991A073236E81CC8FBA073236E81CC8F940A4A4C4B24B6B15F2B";
    attribute INIT_1C of inst : label is "400437449734CBB2DD9D01CC8B0399172C0E644DA4D2488200092D844C6E992E";
    attribute INIT_1D of inst : label is "96208006CB61123BA6D99A65C92E5E00E64581CC8B96073226D22B2CC30884B2";
    attribute INIT_1E of inst : label is "56BD37BD7B0730C2236C90019DD1EEDD1EEFD77F40732340E646DD03991F2835";
    attribute INIT_1F of inst : label is "00000000000000000000000000CDF3BDE3498BEF7BCEB137CE739D622FBCE71A";
    attribute INIT_20 of inst : label is "3AB68F4DE59ED47E59F59ED04B3EB1DE1B6FD2D4E800012AAAD50FFAFE602952";
    attribute INIT_21 of inst : label is "5326645719126DB6332B8069C83CB4995B7B6A4916E3DB3B6D9232652D411F34";
    attribute INIT_22 of inst : label is "E365A59161E290E6489915F47E89E4499111023935511196C91544566AAE90B0";
    attribute INIT_23 of inst : label is "0809C4E9FE668C11AA8C06A3677772DD906241A3F1030E4EF01DCA0565034106";
    attribute INIT_24 of inst : label is "319E3880DE2BFC2100402154B274300840020A4D24E8607D52F43E6580102101";
    attribute INIT_25 of inst : label is "6F129905A65161905C651699C5C21821823C4D4D4D4C4C4C0A585B430B607848";
    attribute INIT_26 of inst : label is "FDC2F57DFDF925FD4F51EF05751429964B02F106E192CB6590CB259799641827";
    attribute INIT_27 of inst : label is "BAF26D37AA0931B41BBBF225130484A04DDF91689316A1776BB908773F2F575C";
    attribute INIT_28 of inst : label is "45A24DD994C994CC766D366D370D89448944C722D162D170C994C89A10019519";
    attribute INIT_29 of inst : label is "4C4249A463B34A9B274C12004B0C395261C764CF551A52A72863D78EC5A2F544";
    attribute INIT_2A of inst : label is "34D34B2966A4C777E592DA4532C7EFB143EFFFDE36EDF7FDAC03E80A9C9C6252";
    attribute INIT_2B of inst : label is "78D7340102FFC6FCBE3D2F3E34D40E5C4CCC36F13CDD2A89CDF8044410232DDB";
    attribute INIT_2C of inst : label is "32271B19128D88890825702454E614721978001F15FF96FBC8FEEE66703CCE74";
    attribute INIT_2D of inst : label is "4CEAAD4CA76CCCB3E8CE42F00000775C264F660B5C3159A5F5913AC895444736";
    attribute INIT_2E of inst : label is "B7A2F01F1CF2D27565965455215CBCD2E0540A4EFEB25E0381F35C315ACC44CC";
    attribute INIT_2F of inst : label is "400000000000000000A5CD27B149EC527B349ECDEEC002C99636499AFAFAFEFF";
    attribute INIT_30 of inst : label is "595803940A5022508D652CA15EC35639CBC47B0D58E7C460BF68DE2D3287EC40";
    attribute INIT_31 of inst : label is "D59FE55CD44A89532A2547371CCD598AE2AA9040404F2497D70466A9C59A1448";
    attribute INIT_32 of inst : label is "40883FA4C82A2BCB26130AF4D1E99268C0ECF99E88F0D4CA5565342F9FFA25AD";
    attribute INIT_33 of inst : label is "0A061201E14209D19D5051EA60741441021D185000008274664450781D052121";
    attribute INIT_34 of inst : label is "3019CB971FFFFB973C30B394E1859CFFE187DC28609EF830FF1E502A184D5794";
    attribute INIT_35 of inst : label is "7200000069A453A000A0CF3C73C427039EFB87BB97DFF5F394D1C86E3119C86E";
    attribute INIT_36 of inst : label is "0B82A888828AA26AC15FF7E002748A69A4000000E722074E821000841D3A440E";
    attribute INIT_37 of inst : label is "EE0986F8074C5F138166A3406F8924D61D6C1D7208FCAD04E035C06BBC944442";
    attribute INIT_38 of inst : label is "7ADE77ADC372DCB737FE69F5225FCC97D54F327C09F037B23D916C8B2A38EA94";
    attribute INIT_39 of inst : label is "578B56CAB5AB8DCA6E137993AFBB97DC00073C34B270636CE0C2C9C819F189E7";
    attribute INIT_3A of inst : label is "B722D424910AAF85156A2115C00004043F10F8BE21E23FAB6FDEB5F42D7516F7";
    attribute INIT_3B of inst : label is "49F689B493E50E9F920200DC04650D0900444441454D49416D61AAAAA0A0089E";
    attribute INIT_3C of inst : label is "00000000034C835BF9B7F76FE69B0B25156AA9453CC51505414A528294A50529";
    attribute INIT_3D of inst : label is "FFF97FE2C03390D7037516AA15EE591C03956628C73B6100276C2006F8074C5F";
    attribute INIT_3E of inst : label is "000000000000000000000000000000000000000007993C057FFF5FFAB00EF011";
    attribute INIT_3F of inst : label is "8000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "BFFFF7B9548B1B86372C6E40DFC233C390F0F04252F48950210C2A2E2E77C91E";
    attribute INIT_01 of inst : label is "522A5F02E0108302DFB58DBF5984B508A926649265712DE79E79EE5F48CFF7B7";
    attribute INIT_02 of inst : label is "CB55ED7A230C552694E58C73C307BE1FBE215738E0001CE3F9E36DC802FFFF48";
    attribute INIT_03 of inst : label is "48C6D96595CF5C4CD1D13563C3331998ECC766385C0986C329898A28863AEFEF";
    attribute INIT_04 of inst : label is "A72EB33DCB8AEFFD2EABFF0BAEFF52EBBFD4FB64FDDB333BB33BB33BB3E326DC";
    attribute INIT_05 of inst : label is "F24CF58FBFA76976B57335CE67B304F67DB4CD39A33462FFFBF5BCC8C4B638F1";
    attribute INIT_06 of inst : label is "551155151041154399A49E619DB493D92496DDC3AD36592A44A0EE8B89B7338D";
    attribute INIT_07 of inst : label is "9259659659649651441451441007368BFCDA2FE36ABB20DB8D933FB59F728455";
    attribute INIT_08 of inst : label is "3ED6DBD787CA08263992DB2CD8E54925B8800001C99681B910A5A5A5A5624925";
    attribute INIT_09 of inst : label is "5DC0956DE36504C7B0DF99C96C92494449A598C6E3E4EB2C47CF61865DDE2FFB";
    attribute INIT_0A of inst : label is "A34DB0E1D6189972525B99C043CCEBDED6DF2AAAAAAAAA3CE6CED7096C964A08";
    attribute INIT_0B of inst : label is "BA8E23A50C4EC5CF060E6CE59EBEFA74F7672C70F74387BB3961839A0C1CD9CB";
    attribute INIT_0C of inst : label is "6474661B4E4CC32B21999BBD918C8E8EC269CD18656637392962694BA72BC2EB";
    attribute INIT_0D of inst : label is "D1C75513B471D18C63BB377BA26474641B4F68E3AB231DA71D58C98ECCDDEECC";
    attribute INIT_0E of inst : label is "C5D6B5E7345CE39C6F39CD356D5B56D5E736E482636DD712E3918AF23A3A099E";
    attribute INIT_0F of inst : label is "8000000000000000000000000000000000000000000000000FFFFFFFB12DB696";
    attribute INIT_10 of inst : label is "B4C98CD18645C6A141E55E0781E4E6C2D85B0B0D9675B5B75E63996DB89B1A0D";
    attribute INIT_11 of inst : label is "571DA38E8B8D6E269D1D91DA38E8B8ED1C745C6B7134CD8CD18645C6A758DB7B";
    attribute INIT_12 of inst : label is "ECE3CD132657C366330AAAA82ABCB4D9A2B06281265CB0FA2B8269D1D31DA71D";
    attribute INIT_13 of inst : label is "07B9982ECAD26D31741D0765CC71036DEB9DFB8C669A1B90D2D252525050D0D0";
    attribute INIT_14 of inst : label is "BA76346C6CDDDBBBA76346C9F64CDD9D1B1A3736EEEDD9D1B1A6B3260E0783E6";
    attribute INIT_15 of inst : label is "7237C799A266CD1157F67197738CBB9C65CCE3AE5FEDE420600321312FBCEDD3";
    attribute INIT_16 of inst : label is "BE0C9D899F06B95DAEF8B5CAEC77C7BF9EC26611DCB06ECC8EE5CA6DEECEEE36";
    attribute INIT_17 of inst : label is "1C0E1D87038761E0F1D8783C74FB9CB1F359E766387638763C763C74F6722663";
    attribute INIT_18 of inst : label is "18A2B9D761084200507060D284344082141C1990187299B633A20E46665C8FA6";
    attribute INIT_19 of inst : label is "D4C94DBD637376767B346A5D626F61954BEAA17D619D98760F81F164AF43E07C";
    attribute INIT_1A of inst : label is "C84ECA4ED49D90AC6EE77FF73276924936667919D9B68675975F10F8BCA55D89";
    attribute INIT_1B of inst : label is "8AEF997C5EC67441C8CCCB8633A22E1C8CCC38633A20C323731CC18C58C72C4E";
    attribute INIT_1C of inst : label is "8ECF233A398577CDBE6F723336C674499B9199B6191C62186766DA19DE466473";
    attribute INIT_1D of inst : label is "18C71D99A4C767919D9CC2BBF6DFA7319D13723334CD8CE89B0CCE310C33B369";
    attribute INIT_1E of inst : label is "171E3BDEE747638ECCD3433B48CCCE6179FA6FD39C8CCDB19D1266E46669C767";
    attribute INIT_1F of inst : label is "4000000000000000000000000110CDE62D722193CC52C4632798A588C66F314B";
    attribute INIT_20 of inst : label is "DEEC93D76622C8D270C622C80E18C45D13CB1846648C019154DDEF56D56CADDB";
    attribute INIT_21 of inst : label is "1B8ED239099F9245545551239C79C6C0E05C0F36FB4AE01C56DB77D331040E64";
    attribute INIT_22 of inst : label is "6B82324B90F8CC7719F48E2AAE3DA0C099DDF23181999DC56D9777630334CA64";
    attribute INIT_23 of inst : label is "584C4EB3000E6914AEBBADD44FEB80DE481A38A3F903042A39BD466D4317438E";
    attribute INIT_24 of inst : label is "70963DA89A3FFC4290E55ACCB3777410A42B14A936EEE8C532F8E07960B8AB41";
    attribute INIT_25 of inst : label is "D068361A2914C36124D36CA6D268B2CA28B4E77EE7F66EE72D917FCE2FF9D97E";
    attribute INIT_26 of inst : label is "7DA77631FD9835FC6F1599253145DB692409245AB36D269361B49369369120D1";
    attribute INIT_27 of inst : label is "1C28D1ECBB34CB46361D28D1EC1A5A35B0ED46CF4C6CD6838E944A4713AF674C";
    attribute INIT_28 of inst : label is "1B3DB17367A367A61CD1ECD1ED87347B347B65CD9E8D9E997367A6060CCB6634";
    attribute INIT_29 of inst : label is "72606D36ABC1F966D4F14CCFCB70AE76AED99395E2A362B5DAABE2739B3D177B";
    attribute INIT_2A of inst : label is "326A2B3D34A6C19F814A41110A24C0CF01EBCE2A30080C211809F0E048DC1323";
    attribute INIT_2B of inst : label is "719C3144615540F93E3BB9BC2DB58A576E13321B469D63DD69000504403321D8";
    attribute INIT_2C of inst : label is "F7465DF3AA2EFDD0314670B49F68A67208599B3791FF16F580F443CFDA4793D9";
    attribute INIT_2D of inst : label is "E6BAF4E8F7F8CDE3EA8B74FAAAAAD7FFA7F7FDECC6085EB4CFBA379D13EE843B";
    attribute INIT_2E of inst : label is "DFDBFB9F16FFF45DB7FFFB6EFFDBFF9B8659DECBFEFFFF2035F4C6085A6666EE";
    attribute INIT_2F of inst : label is "8000000000000000033767FBF9FEFEFFBF9FEFEF7FE002F4E7B771DFAAFFABBA";
    attribute INIT_30 of inst : label is "92E8B78EDA314A388D4949654035D65F518000D7597D80693F4E03A1AAA1BC00";
    attribute INIT_31 of inst : label is "AE8BE3F4664CD9B9332667199C04C88636A29AE8CAE1202FD7042154031626FE";
    attribute INIT_32 of inst : label is "083001203B6E022301C0C6840D089006C81070038045D0423F63AA6B81082FF7";
    attribute INIT_33 of inst : label is "B5FBEFFFFD69362EEA8F5A159F8BFC623162E7A800004D8B98C44007E2FAA121";
    attribute INIT_34 of inst : label is "2011366C1041226C13CF6E6F9E7B73249E7913F79E6083CF005F96D16FBAAFE5";
    attribute INIT_35 of inst : label is "DC000000B6D82C5890010413C103FCEF659679626CB28B2E6FBF365820973648";
    attribute INIT_36 of inst : label is "8B8080A0A81778DDF57D5542408B05B6D8000001BDC118B16020800822C5823B";
    attribute INIT_37 of inst : label is "0A0E08FC035239164820E7240FF24254A15CD1F92400FC92E4D1C583D08DDDD8";
    attribute INIT_38 of inst : label is "5C1745E1585415058500C14A08504254212BC17E51F815862C9161AB42BE8860";
    attribute INIT_39 of inst : label is "D7B75E38FAA381E8AE657A4B9C3F8E1C011A3AC0A0758140EB0281E045D0F578";
    attribute INIT_3A of inst : label is "2D061C61000054020AB4010E45862040E1E00F43C00038002E2B970941CB40F1";
    attribute INIT_3B of inst : label is "4B070000060FE120760408FC414F4A4C020005414745454D4848FFFFF0FAAE23";
    attribute INIT_3C of inst : label is "0000000033093455FAABF157EC180BA51128894460055455544A52A894A55129";
    attribute INIT_3D of inst : label is "4001602A800B9D570517128E700A491438152AA8E0AEF1A055DE3408FC035039";
    attribute INIT_3E of inst : label is "000000000000000000000000000000000000000007A0BC0577F97FF8EFF0BFF1";
    attribute INIT_3F of inst : label is "5000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "72323239548B9DD73B8E7740CA0203FC00FF005A44EB8955010448C8C9D6584E";
    attribute INIT_01 of inst : label is "3A0674104A121D42DFB1AD965AACB508A937679EECA924C71C71DDCACCDA7A7A";
    attribute INIT_02 of inst : label is "DF306E1BF586C57610FAF65A7595255D25450FDEE2220909C15434F8A941A360";
    attribute INIT_03 of inst : label is "6042CB24955445C8919125BCB111888C4462232A0A03577961A5A2A22E1ED7EA";
    attribute INIT_04 of inst : label is "262492E50B0CB3B54F2CED53CB3B44F2CED13B24A82A2A2AAA22AAA2A2AD24EF";
    attribute INIT_05 of inst : label is "B26A88B525412512653366B606AD08D5B4D55148290526FBCDF4940E499230C1";
    attribute INIT_06 of inst : label is "DDDD999DDE799F7D6924F4A0393CB6D9249ED94B927AAF2D4672FF13EDFF628F";
    attribute INIT_07 of inst : label is "040000000000000000000000003E17C93C5F24F17E93F8438ED1083C807C66DD";
    attribute INIT_08 of inst : label is "B6D64E83E699303A80324B399B456DABDC008888E5CF01951AA5252525441040";
    attribute INIT_09 of inst : label is "68C011ED40C60750741B5AD9249249C469273CFB40765155A0CD3ABACA863FFD";
    attribute INIT_0A of inst : label is "779FF0BEB318D92E5259DDA6E5F447C6DED27F9F9F9FBEE56ECEDA0124925D77";
    attribute INIT_0B of inst : label is "5CF735E48DA562BD8B15E8BEE3856E1C2B45F71C2B70E15A2FB8C15B060AD17D";
    attribute INIT_0C of inst : label is "6C76641B66ECC323A199DFBFB1ED8ECE8368DD986462A2968945044A068EDB73";
    attribute INIT_0D of inst : label is "D9864713766191CDC333BF7F636C76661B46ECC323231BB6195CD90CCEF5BDCD";
    attribute INIT_0E of inst : label is "1296B02B740C7D8EF794B2DAB2ADAB2AF3755C82722F93156971A3A63B33098D";
    attribute INIT_0F of inst : label is "4000000000000000000000000000000000000000000000000924924926D24922";
    attribute INIT_10 of inst : label is "34CD8DD98646C42F55755755C17EEEEBDD7BADEDB26FBED2B72D4B6494DF7E09";
    attribute INIT_11 of inst : label is "5B1BB30C8D885E369D9991BB30C8D8DD98646C42D1B4CD8DD98646C42FB8493B";
    attribute INIT_12 of inst : label is "5D428BB2BAC2C624A2822222802B749D7650B31ABE8516562AA369D9931BB619";
    attribute INIT_13 of inst : label is "0571703FDFD34DB83E4F83C0F63BD925CD68510945D85982C2C2C2C2C0C04040";
    attribute INIT_14 of inst : label is "6AD6D7AFAB5A54B4A96952D91C7555B56BEBD6D52D2A5A54B4A9F2BACACCB12C";
    attribute INIT_15 of inst : label is "8ECF7979F3C58B15A59A3CE391E71C8F38E479476925A6D656F3521DD01520A9";
    attribute INIT_16 of inst : label is "53ECBAEFE9EBD5EAF54FDEAF56AA7E9EBF5B2EDA975E3E47D4BABB4936A8888B";
    attribute INIT_17 of inst : label is "CDA68E3369A38CDA68E3369A3E8D4BF7126CCA48AB38AB38AB38AB3F9EEBAFB5";
    attribute INIT_18 of inst : label is "FB103D927FF7BF38AE6F6CD2E3344ECC2B9BDB9C2E3AFBBB2777C66FEFEB5F80";
    attribute INIT_19 of inst : label is "CECF871D2B3F6E02693A43ABA82F73C8B53336A6E9DD9EB594F29EEC0F653CA7";
    attribute INIT_1A of inst : label is "C984C984D70993FCA223B3333364926DA4773E1DD9F58664B5C9F74FDDDEBFBF";
    attribute INIT_1B of inst : label is "7AC4B2A5EC64EEFC89D9B57237E6D5CCDFDFD7237E6F77A93D6D4AB4AA5B5584";
    attribute INIT_1C of inst : label is "8ECD6F3E3AFD725DD2D622766E64EEFEF99BFBFBBD4E6E3866779F1DDEDE7E7D";
    attribute INIT_1D of inst : label is "9B8E19DDF5C767B79F1F7EB12CA97B91BF3622766D78C9DDF5DEA7371C333BCB";
    attribute INIT_1E of inst : label is "6B2F1ADEA7E2C70CEEFAC3335BCDCEBF5C9774B5CCDFDF91BF37BE44ECDEEF53";
    attribute INIT_1F of inst : label is "40000000000000000000000003B8D967A9AF71B2CF535EC3659EA6BD86EB3D4D";
    attribute INIT_20 of inst : label is "E258DC42EAE3DDD27B52E3DC8F2A5C7F81ED4B64E70644AAAA0C95FE7FA4C5CB";
    attribute INIT_21 of inst : label is "35B4922FA08900054551410368117B50AA15413E3B68AA17DB6DA1931C4515C6";
    attribute INIT_22 of inst : label is "5EA25656BB78CC6F6C6483A2A3C9210308CC9160ACCCCD5DB6E2222551115660";
    attribute INIT_23 of inst : label is "D808340BFE9091FB145551144CCDB0CE48181883E9C3022278AC402900158503";
    attribute INIT_24 of inst : label is "419C1D80BBE3B95214C01A9D3BE06454852244A0B7C0C84926280B2E81B03B01";
    attribute INIT_25 of inst : label is "D86C261329948341A6934CA6D36C228A2812BAA223BAA22334B3368866D133B4";
    attribute INIT_26 of inst : label is "3FA33E99EC81937D2546112731C68E49341D269B3A6926DA4124936D249060D1";
    attribute INIT_27 of inst : label is "1B1BD2FF19FFFF4A3F1A9BD2FFFFFA5DF8D4DED7FFED57E3654D58C23284C2C2";
    attribute INIT_28 of inst : label is "FA5FF7AF4FEF4BEEAFD3FFD2FFBBF4FFF4BFEEFDBFFDAFFABF4BFED43CEF4B3D";
    attribute INIT_29 of inst : label is "6A3C2F97A97D51759AAD7CCAA130DF26ACD9D3B0F2F9783BFBA93173BA5F633F";
    attribute INIT_2A of inst : label is "A0EA0D3CD555A7FFD243E051BCCE61EF7E2A61FCB70E56B5D01D57BF7B9B51E1";
    attribute INIT_2B of inst : label is "2DBDB6640244505C1F9F983F0B2441407467B5FE7ECEA888E4D0000100653A8A";
    attribute INIT_2C of inst : label is "6764AEB3BA575DDCA2C3FD998EA963FC287B8E26242FCC4C7C4570EC7F41D87C";
    attribute INIT_2D of inst : label is "A330E72A73D6BB501AB7F59AAAAAFD499494B97887B16D3CEF3B279D93EECEDD";
    attribute INIT_2E of inst : label is "CFC9F9AFC669F4BADF496EBB95B76789EABD5695BDEBB3281888C7B16E2222AA";
    attribute INIT_2F of inst : label is "800000000000000002137A4A5E929724A5C92973197FFD2E5DE72FFEAAFFFBE9";
    attribute INIT_30 of inst : label is "08E515805200280985280C203E00C11705A27A13055C22411F040B8181899A00";
    attribute INIT_31 of inst : label is "2F49E780E59CA394768E533944C4C880348010404264840FCA804444A59EB6E0";
    attribute INIT_32 of inst : label is "019C098451481B432182C0A0CE4142274A5E31C1812540587A07CA21952D0F79";
    attribute INIT_33 of inst : label is "A00DFDFFF680C1D33505A000607402DCC095185000003054650D280015052121";
    attribute INIT_34 of inst : label is "CFE673E5E4104CE5D7DF26E4BEF937493EFA672FBFC103DE005F6A80B7F557DA";
    attribute INIT_35 of inst : label is "1000000010402040100175D7DD7F25E2E8A2FA2CE5148946E4D3718BCE637193";
    attribute INIT_36 of inst : label is "D5DFFD77D8155FD53422A0004008041040000000210100810020780802040202";
    attribute INIT_37 of inst : label is "0ACFEAFC025818122820AF140B80085F01444160A4FCAC52F405C20B91655557";
    attribute INIT_38 of inst : label is "5F1785C14050140505FEC570C95FF017D70BFD7E05F8056CABC5590A883ADA01";
    attribute INIT_39 of inst : label is "95085592A48B85D42E217B0B8CBB865C0500B900E17201C2E40385E001F2D17C";
    attribute INIT_3A of inst : label is "53061C600008040010200000024200000000000000002FC42BDA95F3857072AD";
    attribute INIT_3B of inst : label is "0107E492420FBA6AA40848F4404E40464044480E0A080A08446855555F00585A";
    attribute INIT_3C of inst : label is "000000003067B78000000600041BB00C5062831420C00154550000AA00015400";
    attribute INIT_3D of inst : label is "60154002C02283150B550F2A48AA3C544154F8284A2A146655428CCAFC025818";
    attribute INIT_3E of inst : label is "000000000000000000000000000000000000000007B0ABF958055002B00AA005";
    attribute INIT_3F of inst : label is "1000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "363636319115846919D611970AB57C001F00000EC3E200A15A53C02C2D440D07";
    attribute INIT_01 of inst : label is "42D5461A8751505280C9280D9420285506181201810FEDBEF965B0D88CB63636";
    attribute INIT_02 of inst : label is "017603608C59E83550C82824921249124917BC9102856088896C061400C16286";
    attribute INIT_03 of inst : label is "0C808240011451332526CE052333199AEED7764690001112052122B760A53063";
    attribute INIT_04 of inst : label is "D9A30542161140241050090414024105009002002088088088808800888A0902";
    attribute INIT_05 of inst : label is "20002A2A8ACED96D8718D860221A0443201330C0180303498203609607FE31F4";
    attribute INIT_06 of inst : label is "000000040504001450490A41A6CB2490400336805209C2C0348A94024126DB09";
    attribute INIT_07 of inst : label is "000000000000000000000000000113AB344E2CD138B350C36D63003D81604040";
    attribute INIT_08 of inst : label is "080DB1064908AA8999A402429288301000A8A0A073F2899A0D08080809100000";
    attribute INIT_09 of inst : label is "108080328315513324D2129200240016964852108342384346840C31C701A002";
    attribute INIT_0A of inst : label is "4B0D87042699110956DB5110038A8003232C00202020200DDB2B240E01203F75";
    attribute INIT_0B of inst : label is "05A16844098CD18D56AC7B04268C6AB563D8213063458B1EC109A31AAD58F608";
    attribute INIT_0C of inst : label is "4949420024928032801126332149292A400492500650D984E9D1974E24AB0616";
    attribute INIT_0D of inst : label is "250064524940190900224E764249494200249280328A924801D494008939D90A";
    attribute INIT_0E of inst : label is "41718C6ED2501602448C28A2ECBB2E8A90081240E46F160048442AC0A4A10409";
    attribute INIT_0F of inst : label is "8000000000000000000000000000000000000000000000000492492490092490";
    attribute INIT_10 of inst : label is "4920092500650846F81AC1B078119192324648400C4E9340CCD874DA07127106";
    attribute INIT_11 of inst : label is "D4124A00CA108D0922542324A00CA0925006508448492009250065084440DB62";
    attribute INIT_12 of inst : label is "C484006A099E80A8C077D7D77F8283224AA84BB409830EC46670922548324801";
    attribute INIT_13 of inst : label is "08C88849480C924609C270982860336D8850AA91803E7AB3F1F3F1F3F3F1F3F1";
    attribute INIT_14 of inst : label is "79F1F1E1E3C3C7878F0F1E114413DC7CF878F0F1E1E3C3C7878A220990A2288A";
    attribute INIT_15 of inst : label is "EBEA1A464C9932643A460820B0410582082C10411B6DC1486342E6241FE36C30";
    attribute INIT_16 of inst : label is "50BAEA9CA856351A8D4231A8D56A15BD901B64D99B8576EECCDC26DBEDDDDEEA";
    attribute INIT_17 of inst : label is "D96CC2B65B30AD96CC2B65B308804292288D809A440A440A440A440B0BAA72AB";
    attribute INIT_18 of inst : label is "A78205102D4350B28FCE4E4DB593662CA3F392D8EB2826CC400048800082EEA2";
    attribute INIT_19 of inst : label is "6CC4A4316709F238220A8C06186D5208B1311E2798156F10C438879881610C21";
    attribute INIT_1A of inst : label is "6C806C806D00D881777777762C9B6D9249422E0156D0414539C87643140022A4";
    attribute INIT_1B of inst : label is "7CE43B218AAA122D542450F5401143D542450745080434920850AC2A82156380";
    attribute INIT_1C of inst : label is "008C0743083E621910C544000488000C32200031A4824920054948015C0E8610";
    attribute INIT_1D of inst : label is "9248015250004603A1061F310C8872AA008A55091619542458D241249002A4A0";
    attribute INIT_1E of inst : label is "D3EF9B9EE7002400A92820A381D2C30F9C876439554245A284020E8800086920";
    attribute INIT_1F of inst : label is "40000000000000000000000000689110E618D12221CC31A24443986344A88730";
    attribute INIT_20 of inst : label is "6E36EDD1808BB46C58308BB41B0611728168C204E92100440019A5545520058B";
    attribute INIT_21 of inst : label is "B328669689986DB40011100A5025B902D84B02DA0CB2D85B0DA440662C501137";
    attribute INIT_22 of inst : label is "9B69A59978E69D665019A5AA20B048D09999E11939999990D266667673359500";
    attribute INIT_23 of inst : label is "4008A851040140414141140006651A8C0141451020106F74F696A9A5B41A2204";
    attribute INIT_24 of inst : label is "43980C019B86B410043010CCFB2754061185063AB64EA844CC29616460800801";
    attribute INIT_25 of inst : label is "000002012090412092482110080006182002666667666666227FED89FDB13FEC";
    attribute INIT_26 of inst : label is "02630904B085380370D42608451478000204B04C20200249209248018001106D";
    attribute INIT_27 of inst : label is "9282201055930080489202201089840E44901140B014191263414B30AA00B0B8";
    attribute INIT_28 of inst : label is "8C06490884508051422110201040884408041422910281050880591842A8814A";
    attribute INIT_29 of inst : label is "65372D13EB3161592301408A89000B42E8CC6494D29922056BEB50188C068AA0";
    attribute INIT_2A of inst : label is "0848800824501C404040A860434E0E1EC18B290A256AAD6BA02154C12C482999";
    attribute INIT_2B of inst : label is "0A5B256684414705C04508326FB71B765208271580A88954204D100402800E46";
    attribute INIT_2C of inst : label is "1473860AB1C10119C6C637B79CAB66342A5FAE3706802804081DD0C054898C44";
    attribute INIT_2D of inst : label is "6630C02930BE0AF816032C80000022201DB494D986E1423330AB18518C0AE384";
    attribute INIT_2E of inst : label is "D85B0BC026196C1996D96208B1D2E619471CCD8300DB7343D009C6E140666666";
    attribute INIT_2F of inst : label is "0000000000000000013266DA49B6926DA49B69273920010A13830ACD55000100";
    attribute INIT_30 of inst : label is "6E43D2D34B41A3412438963AFFACA1C4B5357CA28612B55F10B52B13D9551360";
    attribute INIT_31 of inst : label is "64081502B43786D0DA1B40AD02E9952B52C284040401568028A354CF3963C640";
    attribute INIT_32 of inst : label is "7EB0A356ED282F1AB64B288AF005AB781FDF75EBAD2CA6A550150670531F3423";
    attribute INIT_33 of inst : label is "8A161201E8A40E2DDAF2280B9F8BFDAA844AE7A80001032B93F208004AFAA121";
    attribute INIT_34 of inst : label is "281473E4038E00E437DF26E4BEF937003EF8072FBEFFFFDFFFDE222C584AAF88";
    attribute INIT_35 of inst : label is "000000000000000000010C37830725F2E082F820E4107106E493724829937250";
    attribute INIT_36 of inst : label is "FD5D75D7581FFF5575F777600000000000000000000000000000500000000000";
    attribute INIT_37 of inst : label is "01E00A1DC4036101A54A0852A07367231428041A93FF014812240448240FFD55";
    attribute INIT_38 of inst : label is "806018060180601810FF2036000F8603C000012ED4BB504002201000000002A4";
    attribute INIT_39 of inst : label is "003C01200300702380040060300018000484062404044A080890100800030201";
    attribute INIT_3A of inst : label is "9E8E38E000000000000001044240000000000000000007C601C100FCE0360008";
    attribute INIT_3B of inst : label is "B2AC1249255FFF4CC61001B400050006010E0001030301010541AAAAF0AAF7DC";
    attribute INIT_3C of inst : label is "000000003C000820044008800AB44452AA9554AA55F2AAA9AAB5AD556B5AAAD6";
    attribute INIT_3D of inst : label is "201000004020020008C0080024802200470080008600050F5000A1EA1DC40961";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000001200000804000010080000";
    attribute INIT_3F of inst : label is "C800000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "24242426C225AECB4C9299C03D266000000000D94A0C2BE5130035D151660B8F";
    attribute INIT_01 of inst : label is "6760EE079650964DC8DB292003210C2784D55B6D555A4934D34D2B01B6942424";
    attribute INIT_02 of inst : label is "20D5372D9CC38C3050996B0D32C0D300D3042588EFE82265EFFC7C1354C1E399";
    attribute INIT_03 of inst : label is "899249249095491225244C0823331112CCD4441614828192412126466A8D9057";
    attribute INIT_04 of inst : label is "5CA4934001104024841009200002480000920124AA00800088880000884A49B7";
    attribute INIT_05 of inst : label is "9272232FBF87F87F9B9ADD60201A4403241114E69CD39904900800A7342442D6";
    attribute INIT_06 of inst : label is "00000004400400065249E948925992492491339CE45DB6E83592B822F096CB24";
    attribute INIT_07 of inst : label is "0000000000000000000000000018B6B826DAE09B698242026828002000A5D144";
    attribute INIT_08 of inst : label is "0900012E452220C988924922B29D225C12A8AA007CA80903098D8D8D8C000000";
    attribute INIT_09 of inst : label is "13888037911419316449524924924914964C52949139965B42400B2DB330A480";
    attribute INIT_0A of inst : label is "CB299ACB6618325AE4C8728019999821313CAACACACACB35492B7489249262AA";
    attribute INIT_0B of inst : label is "2D2B4AC8590C812904094ECB640948204A765B244A512253B2D9225289129D96";
    attribute INIT_0C of inst : label is "5B5B5927ACB698748C366D2B214B6B6924F196D30E8588ACEB58975AD4AB24B4";
    attribute INIT_0D of inst : label is "6D30E8D25B4C3A4B186CDA56425B5B59278CB698741A12DCC3E0B061B3611948";
    attribute INIT_0E of inst : label is "0139C82A59329252D4A569A6E9BA6ADB999DB364E30020644AC52AC9ADAC93D9";
    attribute INIT_0F of inst : label is "8000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "DBB3C96D30E9668840B10B42C0B3B3B676CEDADA644A4105804AD2012C2A4893";
    attribute INIT_11 of inst : label is "E592DA61D2CD101B76D6792DA61D2C96D30E966880DBB3C96D30E9668A4C924C";
    attribute INIT_12 of inst : label is "E6B3326AC99789A68C82A8022A969976CBA44AF4C991E40CA321B76D67B2DCC3";
    attribute INIT_13 of inst : label is "262644A92A64B26C5B56D5B56966424932D3A64D19381EC2C2C0C0C2C2C2C0C0";
    attribute INIT_14 of inst : label is "D0A4A149429285250A4A1492009349285250A4A14942928525080449A5BB6CD9";
    attribute INIT_15 of inst : label is "0A0A90464C99326461241B6DA0DB6D06DB6836DB924889D946CAC6C4F44B9562";
    attribute INIT_16 of inst : label is "54D6D2952A54A552A952A52A954A912D00934099332544A8C99924922911100A";
    attribute INIT_17 of inst : label is "4160B650582D94160B650582D902D61C25D835B936D936D936D936DA954A54AA";
    attribute INIT_18 of inst : label is "0608C76194200020B848482FC00B68082E1212D4AAAD264C8E4C891C99568E51";
    attribute INIT_19 of inst : label is "24C424A22B4CE310000160F3CA499C310162282D1C326C0B0520A51E30814829";
    attribute INIT_1A of inst : label is "6D436D437E86DAA64444444444DB6DB6DB4B244326CB30D8A10A4252B20022D0";
    attribute INIT_1B of inst : label is "D0A529295991C991239322C48E4CAB1239322C58E5DA981C5AD2956956B48943";
    attribute INIT_1C of inst : label is "61B22B8515684290148CD9EDDAB3DBB16ACF6ED4C0D659C30C9B24C324570822";
    attribute INIT_1D of inst : label is "9670C326CB30D815C20AB4294A4A466CF6EC59EDDAB167B762606B2CE1864D96";
    attribute INIT_1E of inst : label is "D52A495AD31038619365986C8AE1045A14A5252B367B7624F6645891C9953035";
    attribute INIT_1F of inst : label is "80000000000000000000000000E59635F759CB2C6BEEB39658D7DD672C91AFBA";
    attribute INIT_20 of inst : label is "66B68CF5959A9626CC959A9789D2B352E13A564570090111546EA957556A21C3";
    attribute INIT_21 of inst : label is "B7296FA60DD86C96232ABCA6522530369ED3C2D94DD61EC32480486ECEF2A934";
    attribute INIT_22 of inst : label is "EC78849660A69F6E521BE9FC7CB27870BBDDE41427FDDF12405FF76C4BBD189B";
    attribute INIT_23 of inst : label is "610DE9FEFBFAECEFFFABABE95EF7328C9270610422064E666DF4C97D24370A44";
    attribute INIT_24 of inst : label is "84988E02AB0232CE77A7AD85B103C8B18D69EB6A1407918DB29AF21D62C22C05";
    attribute INIT_25 of inst : label is "6CB6592CB65B2492CF67B3D9ECF24F2CB2E644444555555442D8493109221849";
    attribute INIT_26 of inst : label is "42EB4BAC3711688352D99844653428924926592C2D96D92492DB6492C924896D";
    attribute INIT_27 of inst : label is "53026F33994A89BD1953026F33654DE8CA981339A933A32A5B815C362DCCB6B7";
    attribute INIT_28 of inst : label is "CDE62759B8C9BCCE966E326F33B59B8C9BCCED666326733A59BCD4C631B1BD19";
    attribute INIT_29 of inst : label is "581C29247039669918CEF19763464B4BF1ED62F5DD1A48C96E705B9ACDE67322";
    attribute INIT_2A of inst : label is "C0CC007065C152201B608C30229411B6FECDBD95270E46311903BB0A121440C1";
    attribute INIT_2B of inst : label is "899925D5ABEAA72DC0EE1076BDF0AE1D410426F539AB853210314000000A4C76";
    attribute INIT_2C of inst : label is "0DA9B28654D9432A6C24F42457F614FC3CD89049D5207A2C4A056EE67535C260";
    attribute INIT_2D of inst : label is "44AEB60AA527569D142A0958000057D7FD2D288134A706A19C6D4E36A71971AD";
    attribute INIT_2E of inst : label is "985B0BA074D04951049041802530B592D4D2892A40925AE0240974A702666644";
    attribute INIT_2F of inst : label is "0000000000000000032544969125A44969125A45AA40024C9292488AAAAAABFE";
    attribute INIT_30 of inst : label is "6E90BE92FA437A4221789E2C3F9DA1CEB764FC66863AE4D7003F23B397B19241";
    attribute INIT_31 of inst : label is "492A0624BD76AED5DAB95D2574C999207E9004040409A488399645CFBD7AF794";
    attribute INIT_32 of inst : label is "7EFD3224EBE8732F27738844D899D26C118EFDDF8A3FCCE2624646F213BB8948";
    attribute INIT_33 of inst : label is "35F9EFFFE28B31D66520A3F4607408220B2518500000CC946828807FA5052121";
    attribute INIT_34 of inst : label is "EFF72449F4516E49E38E4C491C72626D9C7372471C40038E005EA0D367BD57A8";
    attribute INIT_35 of inst : label is "0000000000000000002079E39E7E48F44D34734E49A68A6C492627D3EFF627DB";
    attribute INIT_36 of inst : label is "F557D5FD581F5D57FDD7D7C00000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0BEFE2A1C0000012010AA000AA000054014001400000A000A005400A8007D57D";
    attribute INIT_38 of inst : label is "505415054150541505FE0170005F8017C00BFC50C54315822C11608B02A80200";
    attribute INIT_39 of inst : label is "45815608B02AF1400A005002802800140000280404500808A010114001400141";
    attribute INIT_3A of inst : label is "263618600000000000000100000200000000000000002F800BC005F0017000B0";
    attribute INIT_3B of inst : label is "AAAC36DB655AAE70F820019608040004010601010303030307035555055500BA";
    attribute INIT_3C of inst : label is "000000002D7FBFE3FDC7FB8FEAB8007003801C0055F7C00300AD6A015AD402B5";
    attribute INIT_3D of inst : label is "6011602AC0229055004510AA008A4154011502A8022C800F159001E2A1C00800";
    attribute INIT_3E of inst : label is "000000000000000000000000000000000000000005102C055804580AB008B015";
    attribute INIT_3F of inst : label is "C800000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "36363639449A19B4336866469FF1A000000000384E0190B0C8642BEDEDE23939";
    attribute INIT_01 of inst : label is "20682C004F02E13FB3208CB2488CB4688D2EE492EDA36DC71C71DC4A48E63636";
    attribute INIT_02 of inst : label is "DE466D9B75AEA1B706F6D6B9658B965B9672874E1888206AB8C0C4C8518142C8";
    attribute INIT_03 of inst : label is "6442492491C15CE89191A4259999CCCC6663332C5ECBDE4B6D8D9BB3243A6846";
    attribute INIT_04 of inst : label is "3204926421249212492484924921249248492124AAA088880000000088E5240C";
    attribute INIT_05 of inst : label is "9248239AEA800000656322926CB50D969256E308610C25B2CB2492084CB7A089";
    attribute INIT_06 of inst : label is "0000000445044107292434A199341249249ECC4389330D9DE0CCE6038C9FB084";
    attribute INIT_07 of inst : label is "000000000000000000000000002E36A938DAA4E36A93244B8C81093484704040";
    attribute INIT_08 of inst : label is "64B64C87248F862719924938094449338828AAAB2A0000251287070704600000";
    attribute INIT_09 of inst : label is "28C1B0C843C0C4E310C91849249249C24D2308C343244186A65960C3088612CB";
    attribute INIT_0A of inst : label is "2084E1B082C8D9A656DB9919C5C44786CEC22A8A8A8A8A3066C48A1924926AAA";
    attribute INIT_0B of inst : label is "51B46D246C24588462C421B082442112210D84162118B1086C20910844884361";
    attribute INIT_0C of inst : label is "642424103E484322E19990A78D6C84848203C908644A6253A0264D018610D746";
    attribute INIT_0D of inst : label is "9086470B2421916CC333235F1B642424101E4843226059221956C30CCC8D7C29";
    attribute INIT_0E of inst : label is "11D4A483160941294E5A9EFA7E8FA7E9CA604C831E6D93997539C4361212083C";
    attribute INIT_0F of inst : label is "4000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "24482C9086469CA354C14C0314CC4C4188310524B7632C9A13250925D0CD0F0C";
    attribute INIT_11 of inst : label is "5A59210C8D3946648909059210C8D2C9086469CA1324482C9086469CA1B24933";
    attribute INIT_12 of inst : label is "394ECD342740C61CB32800028019E6892058E03E2746185201C6489090792219";
    attribute INIT_13 of inst : label is "1D713034959B4D91A4290A4284B98925CD28D138668341181818181A1A1A1A1A";
    attribute INIT_14 of inst : label is "1B33346468C8D191A3234649034E6CCD991A32346468C8D191A013A75A6699A4";
    attribute INIT_15 of inst : label is "0202CB3122448912ACB6208231041188208C41041B6C744C5A631A32150C828D";
    attribute INIT_16 of inst : label is "1644C0DE0B231188C459188C4622C8B180CB63588CD23446C46696DB05999802";
    attribute INIT_17 of inst : label is "8C060863018218C060863018248529E35A28CA49E821E821E821E82591037831";
    attribute INIT_18 of inst : label is "2857999247BDEF8F096163909EE401E1C258590208329D2377B336EF66291519";
    attribute INIT_19 of inst : label is "869B3299A3725C32C870C20C342E618225644CADA19991A4758EB0A1E65D63AC";
    attribute INIT_1A of inst : label is "8064806484C90178222222233B2492492434B099992486648C6B195859DB8919";
    attribute INIT_1B of inst : label is "061585AC6C6EF666DDECCD1B77B3146DDECC51B77B334723A5294294294A1464";
    attribute INIT_1C of inst : label is "0CC9237196830AC2D636377B316EF66285BBD99A39296618666492199646E125";
    attribute INIT_1D of inst : label is "5986199924866591B8C9418D632B0B1BBD98B77B3342DDECCD1C94B30C333249";
    attribute INIT_1E of inst : label is "298B0C6B1B42C30CCC924332C8DC24A0C2B0B58D8DDECCD3BD11A34CE4428E4A";
    attribute INIT_1F of inst : label is "C000000000000000000000000332C9C628A665938C514CCB2718A299964E3145";
    attribute INIT_20 of inst : label is "9548529A4A614991634A61486C294C290D8D29206E0FB0AAAA5DFAAEABACE5CB";
    attribute INIT_21 of inst : label is "739490581CC9DB600114147B2872C249612C27243219612C9249A19030514CC2";
    attribute INIT_22 of inst : label is "2187334991B840E72864162A06490CD9CCCC903984CCCDC9249333272993CB60";
    attribute INIT_23 of inst : label is "CC10F41155511004440045C48545986A4D998EDBC911B710DC9231269892250E";
    attribute INIT_24 of inst : label is "405F448C03E129631CCD189833006658C73A46203600CC2DEA1AE0260998191A";
    attribute INIT_25 of inst : label is "9048241229148241209048241208A68A288A22222222222339896DC92DBD096E";
    attribute INIT_26 of inst : label is "43824E396CDCB6866BA6712310C2964926190412124924924124924824907090";
    attribute INIT_27 of inst : label is "187D91C99925DE46A418FD91C912F23120C3EC8E5CC8C483047E58E4DA28E4E8";
    attribute INIT_28 of inst : label is "323971A6432647206990C991C80A6432647206990C991C81A6472E1C9CCE46A4";
    attribute INIT_29 of inst : label is "72766EB6A9421966F7B7DEEF9F78B434AED19F0D62E3679692A9626332393337";
    attribute INIT_2A of inst : label is "A03A090CA840719830C218110E08404983832938B09135AD76DDB0F4844E9393";
    attribute INIT_2B of inst : label is "1054B31CE35578BA20798C3DE491FA17AC13B21D02089289CFB400000265200D";
    attribute INIT_2C of inst : label is "E7548D73AA46B9D524523CBC9CBA26302C799B3624503CB64050628A1D05120A";
    attribute INIT_2D of inst : label is "2330DB20B1B846E1160B6C60000002B68DB5B64987910B3C4732239951CC8CDA";
    attribute INIT_2E of inst : label is "D85B0B9036596C5D96D9665DBD96F6D9421C458B42DB7BA0748987910C222222";
    attribute INIT_2F of inst : label is "800000000000000001B276DADDB6B76DADDB6B773B7FFE64CB5B60ED55555402";
    attribute INIT_30 of inst : label is "1B6192624D892189C5647DF960C6D16D49BB831B45B5BBC8909CCB05C185BB80";
    attribute INIT_31 of inst : label is "160A11D640580B01602C0ED03A6446CB124FF62626233B5C3DC5B3650B162F67";
    attribute INIT_32 of inst : label is "0190CDBB39310B6B99C8F0374C7E9DA66B62464A7714A60B9D59902A4D491633";
    attribute INIT_33 of inst : label is "8007FDFFE8A0C7799F8228019FDFE088B09AE7A80000306B862888001AFAA121";
    attribute INIT_34 of inst : label is "EFF776EDF7DF6EEDF7DF6EEDBEFB776DBEFB776FBEFFFFDFFFFE82009FF7FFA0";
    attribute INIT_35 of inst : label is "000000000000000000217DF7DF7F6DF6EDB6FB6EEDB6FB6EEDB777DBEFF777DB";
    attribute INIT_36 of inst : label is "00A880AAA00AA282A002A8000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "A010181E3FFFFC01FEF01FFF01FFFF43F43FF03FF0001FF81FF03FE07FE80282";
    attribute INIT_38 of inst : label is "00000010240902400001F40FFD007F403FA0010F243C907C83E41F20FC87FDFF";
    attribute INIT_39 of inst : label is "907E41F20FC8003F81FC0FE07E07FF03FFFE07FBF80FF7F01FEFE03FF03FF000";
    attribute INIT_3A of inst : label is "4140C308000000000000010000020000000000000000007FA03FD00FF40FFA0F";
    attribute INIT_3B of inst : label is "5AAC36DB65551580FE400195000501050107000200000000050100000000008E";
    attribute INIT_3C of inst : label is "000000000CCD655D54BAA9754ABFFFFFFFFFFFFF557D5555555AD6AAB5AD556B";
    attribute INIT_3D of inst : label is "1FE41FC83FC86F90FF90EF21FF21BE43FE42FC87FC837FF0C06FFE181E3FF7FC";
    attribute INIT_3E of inst : label is "000000000000000000000000000000000000000000EE03F907F907F20FF20FE4";
    attribute INIT_3F of inst : label is "C000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "12121211C0010A8215042AC05FE2A000000000380E055008812221C7C6913829";
    attribute INIT_01 of inst : label is "226868002E02823FB2900D92D90CBC018404400044D124820820884508A21212";
    attribute INIT_02 of inst : label is "5D2680C0402805A6068310A1041A105A10420C6E1A800AE03084C825053E1C28";
    attribute INIT_03 of inst : label is "E0024924918558A1020280051111888C44622370CA594A8925050AA002212004";
    attribute INIT_04 of inst : label is "0404922C6165963059658C165963059658C16124800088888888888800440090";
    attribute INIT_05 of inst : label is "925A0310300490494502175624440488B2DA220440881492DB2496102C922080";
    attribute INIT_06 of inst : label is "00000004451001122000908090009249249A45061B041034804082021C9E1004";
    attribute INIT_07 of inst : label is "000000000000000000000000002D1288944A2251288920314480F69479409100";
    attribute INIT_08 of inst : label is "64964C06240D0C4008924D30010C000390A82222800000070B8D8D8D8C000000";
    attribute INIT_09 of inst : label is "204090A501818801004910492492498000060087012C8208A2484104100C164B";
    attribute INIT_0A of inst : label is "818CD0D142D851D65249111B850007025A500020202020104242580924926AAA";
    attribute INIT_0B of inst : label is "68BA2E846824588C62C460D142C4631623068A1223089118345091184488C1A2";
    attribute INIT_0C of inst : label is "5200000034000222C11100E50D6A400000068000445D516A01052008041853A2";
    attribute INIT_0D of inst : label is "0004468E0001116A822201CA1B5200000034000222D0F0041152A6088807282B";
    attribute INIT_0E of inst : label is "1340070212C18031C46B575C371DC7718954AA411B25508B56A9461500000028";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "928038000446570354A40A0294AA2A21442886AD9343249D33269B6CE9EC2D05";
    attribute INIT_11 of inst : label is "597000088CAE0252500007000088CB8000446570329280380004465703EADB6A";
    attribute INIT_12 of inst : label is "352B440C4010451611000002AA95D2548048401E402228280145250000500411";
    attribute INIT_13 of inst : label is "16A8A8385F4924A9D2749D2740C89B6CAEA0402D220300981818181A1A1A1A1A";
    attribute INIT_14 of inst : label is "8D191830306060C0C1818301018066468C0C181830306060C0C002C05D6F5BD2";
    attribute INIT_15 of inst : label is "02028A2204081022C4B3C1451E0A28F05147828A092610844C220C4225588746";
    attribute INIT_16 of inst : label is "1444C0CE0A231188C451188C46228890C08A3150886234468443124904888802";
    attribute INIT_17 of inst : label is "D82C14360B050D82C14360B05086B5D109702D20B050B050B050B05091033831";
    attribute INIT_18 of inst : label is "2047911006B5AD0C114141028A40034304505086410100804200108400351C88";
    attribute INIT_19 of inst : label is "568A0291A2215A1244207814562541066D4CC5A8811100803506A081E44D41A8";
    attribute INIT_1A of inst : label is "0060006014C001F422222222295249249212A991100004448C2A095061FF8089";
    attribute INIT_1B of inst : label is "861505A87008400610800E9842003A610800E9842001A283D6A1035035A91860";
    attribute INIT_1C of inst : label is "0889222197430A82D4380420030840074C21000D143554104440001116444126";
    attribute INIT_1D of inst : label is "550411100004449110CBA18D436A1C021001842001A61080068A1AAA08222000";
    attribute INIT_1E of inst : label is "ADC38C6B1A01820888000222488865D0C6A195060108004A1088D12A5223450D";
    attribute INIT_1F of inst : label is "8000000000000000000000000202810425D40502084BA80A041097501408212E";
    attribute INIT_20 of inst : label is "4DA4699D0D518543538D5184EA71AA309D4635604607802AAA1172A8AAC4CC99";
    attribute INIT_21 of inst : label is "51104850088949211000146A20228249412822006949412892498148210008A3";
    attribute INIT_22 of inst : label is "6905210910B400E62052142A2C402C588888821B10888C8924C2222221128804";
    attribute INIT_23 of inst : label is "C800D04441551450504405D2844E504924988A83E1029202CC80512008110404";
    attribute INIT_24 of inst : label is "405504C0026121D6B181189821014475AC60462012028829B856C00701903980";
    attribute INIT_25 of inst : label is "00000000201000000000000000018010410C2222222222223089248924910925";
    attribute INIT_26 of inst : label is "400240A120D296802A06D80620A2440002100042000000000000000000015000";
    attribute INIT_27 of inst : label is "1055008166008C020010D500810060100086A804088040020A2A088402080408";
    attribute INIT_28 of inst : label is "201021D40204020075008100801D40204020035008100800D4020416188C0200";
    attribute INIT_29 of inst : label is "33272692A887094216C7D88F9E20B810A8C1020902C1279302A8824220102CC2";
    attribute INIT_2A of inst : label is "906908A480807198114008308E0C20CC02204238A08114A55A14201484029919";
    attribute INIT_2B of inst : label is "0050A31C630030A020608431C001F0032003A20D06090001AE80000000568450";
    attribute INIT_2C of inst : label is "5552142AA90A155564422C9C89DA22220C399A22AC6030A64010619D0D033118";
    attribute INIT_2D of inst : label is "23925B60909A446902092448000028160C9096489392839AA6AA935509AA8A68";
    attribute INIT_2E of inst : label is "48090180120B2448B24B3659948652CB02484489404929E07400939286222222";
    attribute INIT_2F of inst : label is "4000000000000000019632484C92132484C92132113FFE54A959506400000002";
    attribute INIT_30 of inst : label is "9121902240812081414C38BC40431E285E49810C78A149C180184A0502852480";
    attribute INIT_31 of inst : label is "120A089520640C819032040830400A4A30000404040321283146000001020526";
    attribute INIT_32 of inst : label is "01A045A139001A6B09D0D0144C2890A62B2202405714445A0940802A20011212";
    attribute INIT_33 of inst : label is "8A1A1201EA8C0CAEEAAAA20A212A002804600800000103803800000060002121";
    attribute INIT_34 of inst : label is "EFF776EDF7DF6EEDF7DF6EEDBEFB776DBEFB776FBEFFFFDFFFDEA22C684AAFA8";
    attribute INIT_35 of inst : label is "000000000000000000017DF7DF7F6DF6EDB6FB6EEDB6FB6EEDB777DBEFF777DB";
    attribute INIT_36 of inst : label is "AA0000AAA808800A20A800000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "340003400000014400034000340000680280068004004003400A80150018888A";
    attribute INIT_38 of inst : label is "AF2BCAE298A6298ACA00068001A00068003400A002800A005002801400500000";
    attribute INIT_39 of inst : label is "0A002801400502801400A005005000280000500000A0000140000280028002BC";
    attribute INIT_3A of inst : label is "60204000000000000000000000000000000000000000500034001A0006800340";
    attribute INIT_3B of inst : label is "02AFC924955545FF0080009C000C000400040008080808080C0055555555558D";
    attribute INIT_3C of inst : label is "000000001A000000020004000AB0000000000000556000000000000000000000";
    attribute INIT_3D of inst : label is "80068005000D000A001A0014003400280068005000D000000A00000140000001";
    attribute INIT_3E of inst : label is "00000000000000000000000000000000000000000A005000A001A00140034002";
    attribute INIT_3F of inst : label is "1000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
